`timescale 1ps / 1ps
/*****************************************************************************
    Verilog RTL Description
    
    Configured at: 07:05:16 CST (+0800), Friday 26 May 2023
    Configured on: ws26
    Configured by: m111064503 (m111064503)
    
    Created by: Stratus DpOpt 21.05.01 
*******************************************************************************/

module SobelFilter_Add_7U_7_4 (
	in1,
	out1
	); /* architecture "behavioural" */ 
input [6:0] in1;
output [6:0] out1;
wire [6:0] asc001;

assign asc001 = 
	+(in1)
	+(7'B0000001);

assign out1 = asc001;
endmodule

/* CADENCE  urjwTQE= : u9/ySxbfrwZIxEzHVQQV8Q== ** DO NOT EDIT THIS LINE ******/



