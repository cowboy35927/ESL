`timescale 1ps / 1ps
module SobelFilter_DivRem_4(
          in1,
          in2,
          out1,
          clk,
          stall
);
   input [48:0] in1;
   input [23:0] in2;
   output [36:0] out1;
   input clk;
   input stall;
wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13,
     n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25,
     n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37,
     n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49,
     n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61,
     n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73,
     n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85,
     n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97,
     n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108,
     n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119,
     n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130,
     n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141,
     n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152,
     n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163,
     n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174,
     n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185,
     n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196,
     n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207,
     n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218,
     n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229,
     n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240,
     n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251,
     n_252, n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262,
     n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273,
     n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284,
     n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295,
     n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306,
     n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317,
     n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328,
     n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339,
     n_340, n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350,
     n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361,
     n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372,
     n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383,
     n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394,
     n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405,
     n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416,
     n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427,
     n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438,
     n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449,
     n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460,
     n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471,
     n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482,
     n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493,
     n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504,
     n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515,
     n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526,
     n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537,
     n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548,
     n_549, n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559,
     n_560, n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570,
     n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581,
     n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592,
     n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603,
     n_604, n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614,
     n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625,
     n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636,
     n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646, n_647,
     n_648, n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658,
     n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669,
     n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680,
     n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691,
     n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702,
     n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713,
     n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724,
     n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734, n_735,
     n_736, n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_746,
     n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755, n_756, n_757,
     n_758, n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768,
     n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779,
     n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790,
     n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801,
     n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812,
     n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820, n_821, n_822, n_823,
     n_824, n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_834,
     n_835, n_836, n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844, n_845,
     n_846, n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856,
     n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865, n_866, n_867,
     n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876, n_877, n_878,
     n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889,
     n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900,
     n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_910, n_911,
     n_912, n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922,
     n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932, n_933,
     n_934, n_935, n_936, n_937, n_938, n_939, n_940, n_941, n_942, n_943, n_944,
     n_945, n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955,
     n_956, n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966,
     n_967, n_968, n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977,
     n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988,
     n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999,
     n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008,
     n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017,
     n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026,
     n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035,
     n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044,
     n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053,
     n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062,
     n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071,
     n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080,
     n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089,
     n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098,
     n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107,
     n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116,
     n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125,
     n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134,
     n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143,
     n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152,
     n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161,
     n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170,
     n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179,
     n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188,
     n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197,
     n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206,
     n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215,
     n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224,
     n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233,
     n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242,
     n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251,
     n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, sub_217_2_n_0,
     sub_217_2_n_1, sub_217_2_n_2, sub_217_2_n_3, sub_217_2_n_4, sub_217_2_n_5,
     sub_217_2_n_6, sub_217_2_n_7, sub_217_2_n_8, sub_217_2_n_9, sub_217_2_n_10,
     sub_217_2_n_12, sub_217_2_n_13, sub_217_2_n_14, sub_217_2_n_15,
     sub_217_2_n_16, sub_217_2_n_17, sub_217_2_n_18, sub_217_2_n_19,
     sub_217_2_n_21, sub_217_2_n_22, sub_217_2_n_23, sub_217_2_n_24,
     sub_217_2_n_25, sub_236_2_n_0, sub_236_2_n_1, sub_236_2_n_2, sub_236_2_n_3,
     sub_236_2_n_4, sub_236_2_n_5, sub_236_2_n_7, sub_236_2_n_8, sub_236_2_n_9,
     sub_236_2_n_10, sub_236_2_n_11, sub_236_2_n_12, sub_236_2_n_13,
     sub_236_2_n_14, sub_236_2_n_15, sub_236_2_n_16, sub_236_2_n_17,
     sub_236_2_n_18, sub_236_2_n_19, sub_236_2_n_20, sub_236_2_n_22,
     sub_236_2_n_23, sub_236_2_n_24, sub_236_2_n_25, sub_236_2_n_26,
     sub_236_2_n_27, sub_236_2_n_28, sub_236_2_n_29, sub_236_2_n_30,
     sub_255_2_n_0, sub_255_2_n_1, sub_255_2_n_2, sub_255_2_n_3, sub_255_2_n_4,
     sub_255_2_n_5, sub_255_2_n_6, sub_255_2_n_7, sub_255_2_n_8, sub_255_2_n_9,
     sub_255_2_n_11, sub_255_2_n_12, sub_255_2_n_13, sub_255_2_n_14,
     sub_255_2_n_15, sub_255_2_n_16, sub_255_2_n_17, sub_255_2_n_18,
     sub_255_2_n_19, sub_255_2_n_20, sub_255_2_n_21, sub_255_2_n_22,
     sub_255_2_n_23, sub_255_2_n_24, sub_255_2_n_25, sub_255_2_n_26,
     sub_255_2_n_28, sub_255_2_n_29, sub_255_2_n_30, sub_255_2_n_31,
     sub_255_2_n_32, sub_255_2_n_33, sub_255_2_n_35, sub_255_2_n_36,
     sub_255_2_n_37, sub_255_2_n_38, sub_255_2_n_39, sub_255_2_n_40,
     sub_255_2_n_41, sub_274_2_n_0, sub_274_2_n_1, sub_274_2_n_2, sub_274_2_n_4,
     sub_274_2_n_5, sub_274_2_n_6, sub_274_2_n_7, sub_274_2_n_8, sub_274_2_n_9,
     sub_274_2_n_10, sub_274_2_n_11, sub_274_2_n_12, sub_274_2_n_13,
     sub_274_2_n_14, sub_274_2_n_15, sub_274_2_n_16, sub_274_2_n_17,
     sub_274_2_n_18, sub_274_2_n_19, sub_274_2_n_20, sub_274_2_n_21,
     sub_274_2_n_22, sub_274_2_n_23, sub_274_2_n_24, sub_274_2_n_26,
     sub_274_2_n_27, sub_274_2_n_28, sub_274_2_n_29, sub_274_2_n_30,
     sub_274_2_n_31, sub_274_2_n_32, sub_274_2_n_33, sub_274_2_n_35,
     sub_274_2_n_36, sub_274_2_n_37, sub_274_2_n_38, sub_274_2_n_39,
     sub_274_2_n_41, sub_274_2_n_42, sub_293_2_n_0, sub_293_2_n_1, sub_293_2_n_3,
     sub_293_2_n_4, sub_293_2_n_5, sub_293_2_n_6, sub_293_2_n_7, sub_293_2_n_9,
     sub_293_2_n_12, sub_293_2_n_14, sub_293_2_n_15, sub_293_2_n_16,
     sub_293_2_n_17, sub_293_2_n_18, sub_293_2_n_19, sub_293_2_n_20,
     sub_293_2_n_21, sub_293_2_n_22, sub_293_2_n_23, sub_293_2_n_24,
     sub_293_2_n_25, sub_293_2_n_26, sub_293_2_n_27, sub_293_2_n_28,
     sub_293_2_n_29, sub_293_2_n_30, sub_293_2_n_31, sub_293_2_n_32,
     sub_293_2_n_33, sub_293_2_n_34, sub_293_2_n_35, sub_293_2_n_36,
     sub_293_2_n_37, sub_293_2_n_38, sub_293_2_n_39, sub_293_2_n_40,
     sub_293_2_n_41, sub_293_2_n_42, sub_293_2_n_43, sub_293_2_n_44,
     sub_293_2_n_45, sub_293_2_n_46, sub_293_2_n_47, sub_293_2_n_48,
     sub_293_2_n_49, sub_293_2_n_50, sub_312_2_n_1, sub_312_2_n_2, sub_312_2_n_3,
     sub_312_2_n_4, sub_312_2_n_5, sub_312_2_n_6, sub_312_2_n_7, sub_312_2_n_9,
     sub_312_2_n_11, sub_312_2_n_12, sub_312_2_n_13, sub_312_2_n_14,
     sub_312_2_n_15, sub_312_2_n_16, sub_312_2_n_17, sub_312_2_n_18,
     sub_312_2_n_19, sub_312_2_n_20, sub_312_2_n_21, sub_312_2_n_22,
     sub_312_2_n_23, sub_312_2_n_24, sub_312_2_n_25, sub_312_2_n_26,
     sub_312_2_n_27, sub_312_2_n_28, sub_312_2_n_29, sub_312_2_n_31,
     sub_312_2_n_32, sub_312_2_n_33, sub_312_2_n_34, sub_312_2_n_35,
     sub_312_2_n_36, sub_312_2_n_37, sub_312_2_n_38, sub_312_2_n_39,
     sub_312_2_n_40, sub_312_2_n_41, sub_312_2_n_42, sub_312_2_n_43,
     sub_312_2_n_44, sub_312_2_n_45, sub_312_2_n_46, sub_312_2_n_47,
     sub_312_2_n_48, sub_312_2_n_49, sub_312_2_n_50, sub_312_2_n_52,
     sub_312_2_n_53, sub_312_2_n_54, sub_312_2_n_55, sub_312_2_n_56,
     sub_331_2_n_1, sub_331_2_n_2, sub_331_2_n_3, sub_331_2_n_5, sub_331_2_n_6,
     sub_331_2_n_7, sub_331_2_n_8, sub_331_2_n_9, sub_331_2_n_10, sub_331_2_n_12,
     sub_331_2_n_13, sub_331_2_n_14, sub_331_2_n_15, sub_331_2_n_16,
     sub_331_2_n_17, sub_331_2_n_18, sub_331_2_n_19, sub_331_2_n_20,
     sub_331_2_n_21, sub_331_2_n_22, sub_331_2_n_23, sub_331_2_n_24,
     sub_331_2_n_25, sub_331_2_n_27, sub_331_2_n_28, sub_331_2_n_29,
     sub_331_2_n_30, sub_331_2_n_31, sub_331_2_n_32, sub_331_2_n_33,
     sub_331_2_n_34, sub_331_2_n_35, sub_331_2_n_36, sub_331_2_n_37,
     sub_331_2_n_38, sub_331_2_n_39, sub_331_2_n_40, sub_331_2_n_41,
     sub_331_2_n_42, sub_331_2_n_43, sub_331_2_n_44, sub_331_2_n_45,
     sub_331_2_n_46, sub_331_2_n_47, sub_331_2_n_48, sub_331_2_n_49,
     sub_331_2_n_50, sub_331_2_n_51, sub_331_2_n_52, sub_331_2_n_53,
     sub_331_2_n_56, sub_331_2_n_58, sub_350_2_n_0, sub_350_2_n_1, sub_350_2_n_2,
     sub_350_2_n_3, sub_350_2_n_4, sub_350_2_n_5, sub_350_2_n_6, sub_350_2_n_7,
     sub_350_2_n_8, sub_350_2_n_9, sub_350_2_n_10, sub_350_2_n_14,
     sub_350_2_n_15, sub_350_2_n_16, sub_350_2_n_18, sub_350_2_n_19,
     sub_350_2_n_20, sub_350_2_n_21, sub_350_2_n_22, sub_350_2_n_23,
     sub_350_2_n_24, sub_350_2_n_25, sub_350_2_n_26, sub_350_2_n_27,
     sub_350_2_n_28, sub_350_2_n_29, sub_350_2_n_30, sub_350_2_n_31,
     sub_350_2_n_32, sub_350_2_n_33, sub_350_2_n_34, sub_350_2_n_35,
     sub_350_2_n_36, sub_350_2_n_38, sub_350_2_n_39, sub_350_2_n_40,
     sub_350_2_n_41, sub_350_2_n_42, sub_350_2_n_43, sub_350_2_n_44,
     sub_350_2_n_45, sub_350_2_n_46, sub_350_2_n_47, sub_350_2_n_48,
     sub_350_2_n_49, sub_350_2_n_50, sub_350_2_n_51, sub_350_2_n_52,
     sub_350_2_n_53, sub_350_2_n_54, sub_350_2_n_55, sub_350_2_n_56,
     sub_350_2_n_57, sub_350_2_n_58, sub_350_2_n_59, sub_350_2_n_60,
     sub_350_2_n_61, sub_350_2_n_62, sub_350_2_n_63, sub_350_2_n_65,
     sub_350_2_n_66, sub_350_2_n_67, sub_350_2_n_68, sub_350_2_n_69,
     sub_350_2_n_70, sub_350_2_n_71, sub_350_2_n_72, sub_350_2_n_73,
     sub_350_2_n_74, sub_350_2_n_75, sub_350_2_n_76, sub_350_2_n_78,
     sub_350_2_n_79, sub_350_2_n_82, sub_369_2_n_0, sub_369_2_n_1, sub_369_2_n_2,
     sub_369_2_n_3, sub_369_2_n_4, sub_369_2_n_5, sub_369_2_n_6, sub_369_2_n_7,
     sub_369_2_n_8, sub_369_2_n_9, sub_369_2_n_13, sub_369_2_n_15,
     sub_369_2_n_16, sub_369_2_n_17, sub_369_2_n_18, sub_369_2_n_19,
     sub_369_2_n_20, sub_369_2_n_21, sub_369_2_n_22, sub_369_2_n_23,
     sub_369_2_n_24, sub_369_2_n_25, sub_369_2_n_26, sub_369_2_n_27,
     sub_369_2_n_28, sub_369_2_n_29, sub_369_2_n_30, sub_369_2_n_31,
     sub_369_2_n_32, sub_369_2_n_33, sub_369_2_n_34, sub_369_2_n_35,
     sub_369_2_n_36, sub_369_2_n_37, sub_369_2_n_39, sub_369_2_n_40,
     sub_369_2_n_41, sub_369_2_n_42, sub_369_2_n_43, sub_369_2_n_44,
     sub_369_2_n_45, sub_369_2_n_46, sub_369_2_n_47, sub_369_2_n_48,
     sub_369_2_n_49, sub_369_2_n_50, sub_369_2_n_51, sub_369_2_n_52,
     sub_369_2_n_53, sub_369_2_n_54, sub_369_2_n_55, sub_369_2_n_56,
     sub_369_2_n_57, sub_369_2_n_58, sub_369_2_n_59, sub_369_2_n_60,
     sub_369_2_n_61, sub_369_2_n_62, sub_369_2_n_63, sub_369_2_n_64,
     sub_369_2_n_65, sub_369_2_n_67, sub_369_2_n_68, sub_369_2_n_69,
     sub_369_2_n_70, sub_369_2_n_71, sub_369_2_n_72, sub_369_2_n_73,
     sub_369_2_n_74, sub_369_2_n_75, sub_369_2_n_76, sub_369_2_n_78,
     sub_369_2_n_79, sub_369_2_n_80, sub_369_2_n_81, sub_369_2_n_82,
     sub_369_2_n_84, sub_369_2_n_85, sub_369_2_n_86, sub_388_2_n_0,
     sub_388_2_n_1, sub_388_2_n_2, sub_388_2_n_4, sub_388_2_n_5, sub_388_2_n_6,
     sub_388_2_n_7, sub_388_2_n_8, sub_388_2_n_9, sub_388_2_n_10, sub_388_2_n_11,
     sub_388_2_n_12, sub_388_2_n_18, sub_388_2_n_19, sub_388_2_n_20,
     sub_388_2_n_21, sub_388_2_n_23, sub_388_2_n_24, sub_388_2_n_25,
     sub_388_2_n_26, sub_388_2_n_27, sub_388_2_n_28, sub_388_2_n_29,
     sub_388_2_n_30, sub_388_2_n_31, sub_388_2_n_32, sub_388_2_n_33,
     sub_388_2_n_34, sub_388_2_n_35, sub_388_2_n_36, sub_388_2_n_37,
     sub_388_2_n_38, sub_388_2_n_39, sub_388_2_n_40, sub_388_2_n_41,
     sub_388_2_n_42, sub_388_2_n_43, sub_388_2_n_44, sub_388_2_n_46,
     sub_388_2_n_47, sub_388_2_n_48, sub_388_2_n_49, sub_388_2_n_50,
     sub_388_2_n_51, sub_388_2_n_52, sub_388_2_n_53, sub_388_2_n_54,
     sub_388_2_n_55, sub_388_2_n_56, sub_388_2_n_57, sub_388_2_n_58,
     sub_388_2_n_59, sub_388_2_n_60, sub_388_2_n_61, sub_388_2_n_62,
     sub_388_2_n_63, sub_388_2_n_64, sub_388_2_n_65, sub_388_2_n_66,
     sub_388_2_n_67, sub_388_2_n_68, sub_388_2_n_69, sub_388_2_n_70,
     sub_388_2_n_71, sub_388_2_n_72, sub_388_2_n_73, sub_388_2_n_74,
     sub_388_2_n_75, sub_388_2_n_76, sub_388_2_n_77, sub_388_2_n_78,
     sub_388_2_n_79, sub_388_2_n_80, sub_388_2_n_81, sub_388_2_n_82,
     sub_388_2_n_83, sub_388_2_n_84, sub_388_2_n_85, sub_388_2_n_86,
     sub_388_2_n_87, sub_388_2_n_88, sub_388_2_n_89, sub_388_2_n_90,
     sub_388_2_n_91, sub_388_2_n_92, sub_388_2_n_93, sub_388_2_n_94,
     sub_388_2_n_96, sub_388_2_n_97, sub_388_2_n_98, sub_388_2_n_99,
     sub_388_2_n_100, sub_388_2_n_101, sub_388_2_n_102, sub_388_2_n_103,
     sub_388_2_n_104, sub_388_2_n_106, sub_388_2_n_107, sub_388_2_n_108,
     sub_388_2_n_110, sub_407_2_n_0, sub_407_2_n_1, sub_407_2_n_2, sub_407_2_n_3,
     sub_407_2_n_4, sub_407_2_n_5, sub_407_2_n_6, sub_407_2_n_7, sub_407_2_n_8,
     sub_407_2_n_9, sub_407_2_n_10, sub_407_2_n_11, sub_407_2_n_12,
     sub_407_2_n_13, sub_407_2_n_14, sub_407_2_n_15, sub_407_2_n_16,
     sub_407_2_n_17, sub_407_2_n_19, sub_407_2_n_25, sub_407_2_n_27,
     sub_407_2_n_28, sub_407_2_n_29, sub_407_2_n_30, sub_407_2_n_31,
     sub_407_2_n_32, sub_407_2_n_33, sub_407_2_n_34, sub_407_2_n_35,
     sub_407_2_n_36, sub_407_2_n_37, sub_407_2_n_38, sub_407_2_n_39,
     sub_407_2_n_40, sub_407_2_n_41, sub_407_2_n_42, sub_407_2_n_43,
     sub_407_2_n_44, sub_407_2_n_45, sub_407_2_n_47, sub_407_2_n_48,
     sub_407_2_n_49, sub_407_2_n_50, sub_407_2_n_51, sub_407_2_n_52,
     sub_407_2_n_53, sub_407_2_n_54, sub_407_2_n_55, sub_407_2_n_56,
     sub_407_2_n_57, sub_407_2_n_58, sub_407_2_n_59, sub_407_2_n_60,
     sub_407_2_n_61, sub_407_2_n_62, sub_407_2_n_63, sub_407_2_n_64,
     sub_407_2_n_65, sub_407_2_n_66, sub_407_2_n_67, sub_407_2_n_68,
     sub_407_2_n_69, sub_407_2_n_70, sub_407_2_n_71, sub_407_2_n_72,
     sub_407_2_n_74, sub_407_2_n_75, sub_407_2_n_76, sub_407_2_n_77,
     sub_407_2_n_78, sub_407_2_n_79, sub_407_2_n_80, sub_407_2_n_81,
     sub_407_2_n_82, sub_407_2_n_83, sub_407_2_n_84, sub_407_2_n_85,
     sub_407_2_n_86, sub_407_2_n_89, sub_426_2_n_0, sub_426_2_n_1, sub_426_2_n_2,
     sub_426_2_n_3, sub_426_2_n_4, sub_426_2_n_5, sub_426_2_n_6, sub_426_2_n_7,
     sub_426_2_n_8, sub_426_2_n_9, sub_426_2_n_10, sub_426_2_n_11,
     sub_426_2_n_12, sub_426_2_n_13, sub_426_2_n_14, sub_426_2_n_15,
     sub_426_2_n_16, sub_426_2_n_17, sub_426_2_n_22, sub_426_2_n_23,
     sub_426_2_n_25, sub_426_2_n_26, sub_426_2_n_27, sub_426_2_n_28,
     sub_426_2_n_29, sub_426_2_n_30, sub_426_2_n_31, sub_426_2_n_32,
     sub_426_2_n_33, sub_426_2_n_34, sub_426_2_n_35, sub_426_2_n_37,
     sub_426_2_n_38, sub_426_2_n_39, sub_426_2_n_40, sub_426_2_n_41,
     sub_426_2_n_42, sub_426_2_n_43, sub_426_2_n_44, sub_426_2_n_45,
     sub_426_2_n_46, sub_426_2_n_47, sub_426_2_n_48, sub_426_2_n_49,
     sub_426_2_n_50, sub_426_2_n_51, sub_426_2_n_52, sub_426_2_n_53,
     sub_426_2_n_54, sub_426_2_n_55, sub_426_2_n_56, sub_426_2_n_57,
     sub_426_2_n_58, sub_426_2_n_60, sub_426_2_n_61, sub_426_2_n_62,
     sub_426_2_n_63, sub_426_2_n_64, sub_426_2_n_65, sub_426_2_n_66,
     sub_426_2_n_67, sub_426_2_n_68, sub_426_2_n_69, sub_426_2_n_70,
     sub_426_2_n_71, sub_426_2_n_72, sub_426_2_n_73, sub_426_2_n_74,
     sub_426_2_n_75, sub_426_2_n_76, sub_426_2_n_77, sub_426_2_n_78,
     sub_426_2_n_79, sub_426_2_n_80, sub_426_2_n_81, sub_426_2_n_82,
     sub_426_2_n_83, sub_426_2_n_84, sub_426_2_n_85, sub_426_2_n_86,
     sub_426_2_n_87, sub_426_2_n_88, sub_426_2_n_89, sub_426_2_n_90,
     sub_426_2_n_91, sub_426_2_n_93, sub_426_2_n_94, sub_426_2_n_95,
     sub_426_2_n_96, sub_426_2_n_97, sub_426_2_n_98, sub_426_2_n_99,
     sub_426_2_n_100, sub_426_2_n_101, sub_426_2_n_102, sub_426_2_n_103,
     sub_426_2_n_104, sub_426_2_n_105, sub_426_2_n_106, sub_426_2_n_107,
     sub_426_2_n_108, sub_426_2_n_109, sub_426_2_n_110, sub_426_2_n_112,
     sub_426_2_n_113, sub_426_2_n_116, sub_426_2_n_117, sub_426_2_n_120,
     sub_445_2_n_0, sub_445_2_n_1, sub_445_2_n_2, sub_445_2_n_3, sub_445_2_n_4,
     sub_445_2_n_5, sub_445_2_n_6, sub_445_2_n_7, sub_445_2_n_8, sub_445_2_n_9,
     sub_445_2_n_10, sub_445_2_n_11, sub_445_2_n_12, sub_445_2_n_13,
     sub_445_2_n_14, sub_445_2_n_15, sub_445_2_n_16, sub_445_2_n_17,
     sub_445_2_n_19, sub_445_2_n_20, sub_445_2_n_24, sub_445_2_n_25,
     sub_445_2_n_26, sub_445_2_n_28, sub_445_2_n_29, sub_445_2_n_30,
     sub_445_2_n_31, sub_445_2_n_32, sub_445_2_n_34, sub_445_2_n_35,
     sub_445_2_n_36, sub_445_2_n_37, sub_445_2_n_38, sub_445_2_n_39,
     sub_445_2_n_40, sub_445_2_n_41, sub_445_2_n_42, sub_445_2_n_43,
     sub_445_2_n_44, sub_445_2_n_45, sub_445_2_n_46, sub_445_2_n_47,
     sub_445_2_n_48, sub_445_2_n_49, sub_445_2_n_50, sub_445_2_n_51,
     sub_445_2_n_52, sub_445_2_n_53, sub_445_2_n_54, sub_445_2_n_55,
     sub_445_2_n_56, sub_445_2_n_57, sub_445_2_n_58, sub_445_2_n_59,
     sub_445_2_n_60, sub_445_2_n_61, sub_445_2_n_63, sub_445_2_n_64,
     sub_445_2_n_65, sub_445_2_n_66, sub_445_2_n_67, sub_445_2_n_68,
     sub_445_2_n_69, sub_445_2_n_70, sub_445_2_n_71, sub_445_2_n_72,
     sub_445_2_n_73, sub_445_2_n_74, sub_445_2_n_75, sub_445_2_n_76,
     sub_445_2_n_77, sub_445_2_n_78, sub_445_2_n_79, sub_445_2_n_80,
     sub_445_2_n_81, sub_445_2_n_82, sub_445_2_n_83, sub_445_2_n_84,
     sub_445_2_n_85, sub_445_2_n_86, sub_445_2_n_87, sub_445_2_n_88,
     sub_445_2_n_89, sub_445_2_n_90, sub_445_2_n_91, sub_445_2_n_92,
     sub_445_2_n_93, sub_445_2_n_94, sub_445_2_n_95, sub_445_2_n_96,
     sub_445_2_n_97, sub_445_2_n_98, sub_445_2_n_99, sub_445_2_n_100,
     sub_445_2_n_101, sub_445_2_n_102, sub_445_2_n_103, sub_445_2_n_105,
     sub_445_2_n_106, sub_445_2_n_107, sub_445_2_n_108, sub_445_2_n_109,
     sub_445_2_n_110, sub_445_2_n_111, sub_445_2_n_112, sub_445_2_n_113,
     sub_445_2_n_114, sub_445_2_n_115, sub_445_2_n_116, sub_445_2_n_117,
     sub_445_2_n_118, sub_445_2_n_119, sub_445_2_n_120, sub_445_2_n_121,
     sub_445_2_n_122, sub_445_2_n_123, sub_445_2_n_124, sub_445_2_n_126,
     sub_445_2_n_127, sub_445_2_n_128, sub_445_2_n_129, sub_445_2_n_130,
     sub_445_2_n_131, sub_445_2_n_132, sub_445_2_n_133, sub_445_2_n_134,
     sub_445_2_n_136, sub_445_2_n_137, sub_445_2_n_138, sub_445_2_n_140,
     sub_445_2_n_141, sub_445_2_n_143, sub_466_2_n_0, sub_466_2_n_1,
     sub_466_2_n_2, sub_466_2_n_3, sub_466_2_n_4, sub_466_2_n_5, sub_466_2_n_6,
     sub_466_2_n_7, sub_466_2_n_8, sub_466_2_n_9, sub_466_2_n_10, sub_466_2_n_11,
     sub_466_2_n_12, sub_466_2_n_13, sub_466_2_n_14, sub_466_2_n_15,
     sub_466_2_n_16, sub_466_2_n_17, sub_466_2_n_18, sub_466_2_n_19,
     sub_466_2_n_20, sub_466_2_n_21, sub_466_2_n_23, sub_466_2_n_26,
     sub_466_2_n_30, sub_466_2_n_31, sub_466_2_n_33, sub_466_2_n_34,
     sub_466_2_n_35, sub_466_2_n_36, sub_466_2_n_37, sub_466_2_n_38,
     sub_466_2_n_39, sub_466_2_n_41, sub_466_2_n_42, sub_466_2_n_43,
     sub_466_2_n_44, sub_466_2_n_45, sub_466_2_n_46, sub_466_2_n_47,
     sub_466_2_n_48, sub_466_2_n_49, sub_466_2_n_50, sub_466_2_n_51,
     sub_466_2_n_52, sub_466_2_n_53, sub_466_2_n_54, sub_466_2_n_55,
     sub_466_2_n_56, sub_466_2_n_57, sub_466_2_n_58, sub_466_2_n_59,
     sub_466_2_n_60, sub_466_2_n_61, sub_466_2_n_62, sub_466_2_n_63,
     sub_466_2_n_64, sub_466_2_n_65, sub_466_2_n_66, sub_466_2_n_67,
     sub_466_2_n_68, sub_466_2_n_70, sub_466_2_n_71, sub_466_2_n_72,
     sub_466_2_n_73, sub_466_2_n_74, sub_466_2_n_75, sub_466_2_n_76,
     sub_466_2_n_77, sub_466_2_n_78, sub_466_2_n_79, sub_466_2_n_80,
     sub_466_2_n_81, sub_466_2_n_82, sub_466_2_n_83, sub_466_2_n_84,
     sub_466_2_n_85, sub_466_2_n_86, sub_466_2_n_87, sub_466_2_n_88,
     sub_466_2_n_89, sub_466_2_n_90, sub_466_2_n_91, sub_466_2_n_92,
     sub_466_2_n_93, sub_466_2_n_94, sub_466_2_n_95, sub_466_2_n_96,
     sub_466_2_n_97, sub_466_2_n_98, sub_466_2_n_99, sub_466_2_n_100,
     sub_466_2_n_101, sub_466_2_n_102, sub_466_2_n_103, sub_466_2_n_104,
     sub_466_2_n_105, sub_466_2_n_106, sub_466_2_n_107, sub_466_2_n_108,
     sub_466_2_n_110, sub_466_2_n_111, sub_466_2_n_112, sub_466_2_n_113,
     sub_466_2_n_114, sub_466_2_n_115, sub_466_2_n_116, sub_466_2_n_117,
     sub_466_2_n_118, sub_466_2_n_119, sub_466_2_n_120, sub_466_2_n_121,
     sub_466_2_n_122, sub_466_2_n_123, sub_466_2_n_125, sub_466_2_n_126,
     sub_466_2_n_127, sub_466_2_n_128, sub_466_2_n_129, sub_466_2_n_130,
     sub_466_2_n_131, sub_466_2_n_133, sub_466_2_n_134, sub_466_2_n_135,
     sub_466_2_n_136, sub_466_2_n_137, sub_466_2_n_138, sub_466_2_n_139,
     sub_466_2_n_140, sub_466_2_n_141, sub_466_2_n_144, sub_466_2_n_146,
     sub_466_2_n_147, sub_487_2_n_0, sub_487_2_n_1, sub_487_2_n_2, sub_487_2_n_3,
     sub_487_2_n_4, sub_487_2_n_5, sub_487_2_n_6, sub_487_2_n_7, sub_487_2_n_8,
     sub_487_2_n_9, sub_487_2_n_10, sub_487_2_n_11, sub_487_2_n_12,
     sub_487_2_n_13, sub_487_2_n_14, sub_487_2_n_15, sub_487_2_n_16,
     sub_487_2_n_17, sub_487_2_n_18, sub_487_2_n_19, sub_487_2_n_20,
     sub_487_2_n_21, sub_487_2_n_22, sub_487_2_n_23, sub_487_2_n_24,
     sub_487_2_n_29, sub_487_2_n_34, sub_487_2_n_35, sub_487_2_n_37,
     sub_487_2_n_38, sub_487_2_n_40, sub_487_2_n_41, sub_487_2_n_42,
     sub_487_2_n_43, sub_487_2_n_44, sub_487_2_n_45, sub_487_2_n_46,
     sub_487_2_n_47, sub_487_2_n_48, sub_487_2_n_49, sub_487_2_n_50,
     sub_487_2_n_51, sub_487_2_n_52, sub_487_2_n_53, sub_487_2_n_54,
     sub_487_2_n_55, sub_487_2_n_56, sub_487_2_n_57, sub_487_2_n_58,
     sub_487_2_n_60, sub_487_2_n_61, sub_487_2_n_62, sub_487_2_n_63,
     sub_487_2_n_64, sub_487_2_n_65, sub_487_2_n_66, sub_487_2_n_67,
     sub_487_2_n_68, sub_487_2_n_69, sub_487_2_n_70, sub_487_2_n_71,
     sub_487_2_n_72, sub_487_2_n_73, sub_487_2_n_74, sub_487_2_n_75,
     sub_487_2_n_76, sub_487_2_n_77, sub_487_2_n_78, sub_487_2_n_79,
     sub_487_2_n_80, sub_487_2_n_81, sub_487_2_n_82, sub_487_2_n_83,
     sub_487_2_n_84, sub_487_2_n_85, sub_487_2_n_86, sub_487_2_n_87,
     sub_487_2_n_88, sub_487_2_n_89, sub_487_2_n_90, sub_487_2_n_91,
     sub_487_2_n_92, sub_487_2_n_93, sub_487_2_n_94, sub_487_2_n_95,
     sub_487_2_n_96, sub_487_2_n_97, sub_487_2_n_98, sub_487_2_n_99,
     sub_487_2_n_100, sub_487_2_n_101, sub_487_2_n_102, sub_487_2_n_103,
     sub_487_2_n_105, sub_487_2_n_106, sub_487_2_n_107, sub_487_2_n_108,
     sub_487_2_n_109, sub_487_2_n_110, sub_487_2_n_111, sub_487_2_n_112,
     sub_487_2_n_113, sub_487_2_n_114, sub_487_2_n_115, sub_487_2_n_116,
     sub_487_2_n_117, sub_487_2_n_118, sub_487_2_n_119, sub_487_2_n_121,
     sub_487_2_n_122, sub_487_2_n_123, sub_487_2_n_124, sub_487_2_n_125,
     sub_487_2_n_126, sub_487_2_n_127, sub_508_2_n_0, sub_508_2_n_1,
     sub_508_2_n_2, sub_508_2_n_3, sub_508_2_n_4, sub_508_2_n_5, sub_508_2_n_6,
     sub_508_2_n_7, sub_508_2_n_8, sub_508_2_n_9, sub_508_2_n_10, sub_508_2_n_11,
     sub_508_2_n_12, sub_508_2_n_13, sub_508_2_n_14, sub_508_2_n_15,
     sub_508_2_n_16, sub_508_2_n_17, sub_508_2_n_18, sub_508_2_n_19,
     sub_508_2_n_20, sub_508_2_n_21, sub_508_2_n_22, sub_508_2_n_23,
     sub_508_2_n_24, sub_508_2_n_25, sub_508_2_n_26, sub_508_2_n_27,
     sub_508_2_n_28, sub_508_2_n_35, sub_508_2_n_36, sub_508_2_n_37,
     sub_508_2_n_38, sub_508_2_n_39, sub_508_2_n_41, sub_508_2_n_42,
     sub_508_2_n_43, sub_508_2_n_44, sub_508_2_n_46, sub_508_2_n_47,
     sub_508_2_n_48, sub_508_2_n_49, sub_508_2_n_50, sub_508_2_n_51,
     sub_508_2_n_52, sub_508_2_n_53, sub_508_2_n_54, sub_508_2_n_55,
     sub_508_2_n_56, sub_508_2_n_57, sub_508_2_n_58, sub_508_2_n_59,
     sub_508_2_n_60, sub_508_2_n_61, sub_508_2_n_62, sub_508_2_n_63,
     sub_508_2_n_64, sub_508_2_n_65, sub_508_2_n_66, sub_508_2_n_67,
     sub_508_2_n_68, sub_508_2_n_69, sub_508_2_n_70, sub_508_2_n_71,
     sub_508_2_n_72, sub_508_2_n_73, sub_508_2_n_74, sub_508_2_n_75,
     sub_508_2_n_76, sub_508_2_n_77, sub_508_2_n_78, sub_508_2_n_79,
     sub_508_2_n_80, sub_508_2_n_82, sub_508_2_n_83, sub_508_2_n_84,
     sub_508_2_n_85, sub_508_2_n_86, sub_508_2_n_87, sub_508_2_n_88,
     sub_508_2_n_89, sub_508_2_n_90, sub_508_2_n_91, sub_508_2_n_92,
     sub_508_2_n_93, sub_508_2_n_94, sub_508_2_n_95, sub_508_2_n_96,
     sub_508_2_n_97, sub_508_2_n_98, sub_508_2_n_99, sub_508_2_n_100,
     sub_508_2_n_101, sub_508_2_n_102, sub_508_2_n_103, sub_508_2_n_104,
     sub_508_2_n_105, sub_508_2_n_106, sub_508_2_n_107, sub_508_2_n_108,
     sub_508_2_n_109, sub_508_2_n_110, sub_508_2_n_111, sub_508_2_n_112,
     sub_508_2_n_113, sub_508_2_n_114, sub_508_2_n_115, sub_508_2_n_116,
     sub_508_2_n_117, sub_508_2_n_118, sub_508_2_n_119, sub_508_2_n_120,
     sub_508_2_n_122, sub_508_2_n_123, sub_508_2_n_124, sub_508_2_n_125,
     sub_508_2_n_126, sub_508_2_n_127, sub_508_2_n_128, sub_508_2_n_129,
     sub_508_2_n_130, sub_508_2_n_131, sub_508_2_n_132, sub_508_2_n_133,
     sub_508_2_n_134, sub_508_2_n_137, sub_508_2_n_138, sub_508_2_n_139,
     sub_508_2_n_140, sub_508_2_n_141, sub_508_2_n_142, sub_508_2_n_143,
     sub_508_2_n_146, sub_508_2_n_148, sub_508_2_n_149, sub_508_2_n_150,
     sub_508_2_n_151, sub_508_2_n_154, sub_508_2_n_155, sub_529_2_n_0,
     sub_529_2_n_1, sub_529_2_n_2, sub_529_2_n_3, sub_529_2_n_4, sub_529_2_n_5,
     sub_529_2_n_6, sub_529_2_n_7, sub_529_2_n_8, sub_529_2_n_9, sub_529_2_n_10,
     sub_529_2_n_11, sub_529_2_n_12, sub_529_2_n_13, sub_529_2_n_14,
     sub_529_2_n_15, sub_529_2_n_16, sub_529_2_n_17, sub_529_2_n_18,
     sub_529_2_n_19, sub_529_2_n_20, sub_529_2_n_21, sub_529_2_n_22,
     sub_529_2_n_23, sub_529_2_n_24, sub_529_2_n_25, sub_529_2_n_26,
     sub_529_2_n_27, sub_529_2_n_33, sub_529_2_n_41, sub_529_2_n_42,
     sub_529_2_n_43, sub_529_2_n_46, sub_529_2_n_47, sub_529_2_n_48,
     sub_529_2_n_49, sub_529_2_n_50, sub_529_2_n_51, sub_529_2_n_53,
     sub_529_2_n_54, sub_529_2_n_55, sub_529_2_n_56, sub_529_2_n_57,
     sub_529_2_n_58, sub_529_2_n_59, sub_529_2_n_60, sub_529_2_n_61,
     sub_529_2_n_62, sub_529_2_n_63, sub_529_2_n_64, sub_529_2_n_65,
     sub_529_2_n_66, sub_529_2_n_67, sub_529_2_n_68, sub_529_2_n_69,
     sub_529_2_n_70, sub_529_2_n_71, sub_529_2_n_72, sub_529_2_n_73,
     sub_529_2_n_74, sub_529_2_n_75, sub_529_2_n_76, sub_529_2_n_77,
     sub_529_2_n_78, sub_529_2_n_79, sub_529_2_n_81, sub_529_2_n_82,
     sub_529_2_n_83, sub_529_2_n_84, sub_529_2_n_85, sub_529_2_n_86,
     sub_529_2_n_87, sub_529_2_n_88, sub_529_2_n_89, sub_529_2_n_90,
     sub_529_2_n_91, sub_529_2_n_92, sub_529_2_n_93, sub_529_2_n_94,
     sub_529_2_n_95, sub_529_2_n_96, sub_529_2_n_97, sub_529_2_n_98,
     sub_529_2_n_99, sub_529_2_n_100, sub_529_2_n_101, sub_529_2_n_102,
     sub_529_2_n_103, sub_529_2_n_104, sub_529_2_n_105, sub_529_2_n_106,
     sub_529_2_n_107, sub_529_2_n_108, sub_529_2_n_109, sub_529_2_n_110,
     sub_529_2_n_111, sub_529_2_n_112, sub_529_2_n_113, sub_529_2_n_114,
     sub_529_2_n_115, sub_529_2_n_116, sub_529_2_n_117, sub_529_2_n_118,
     sub_529_2_n_119, sub_529_2_n_120, sub_529_2_n_121, sub_529_2_n_122,
     sub_529_2_n_123, sub_529_2_n_124, sub_529_2_n_125, sub_529_2_n_126,
     sub_529_2_n_127, sub_529_2_n_128, sub_529_2_n_129, sub_529_2_n_130,
     sub_529_2_n_132, sub_529_2_n_133, sub_529_2_n_134, sub_529_2_n_135,
     sub_529_2_n_136, sub_529_2_n_137, sub_529_2_n_138, sub_529_2_n_139,
     sub_529_2_n_140, sub_529_2_n_141, sub_529_2_n_142, sub_529_2_n_143,
     sub_529_2_n_144, sub_529_2_n_145, sub_529_2_n_146, sub_529_2_n_147,
     sub_529_2_n_149, sub_529_2_n_150, sub_529_2_n_151, sub_529_2_n_152,
     sub_529_2_n_153, sub_529_2_n_154, sub_529_2_n_155, sub_550_2_n_0,
     sub_550_2_n_1, sub_550_2_n_3, sub_550_2_n_4, sub_550_2_n_5, sub_550_2_n_6,
     sub_550_2_n_7, sub_550_2_n_8, sub_550_2_n_9, sub_550_2_n_10, sub_550_2_n_11,
     sub_550_2_n_12, sub_550_2_n_13, sub_550_2_n_14, sub_550_2_n_15,
     sub_550_2_n_16, sub_550_2_n_17, sub_550_2_n_18, sub_550_2_n_19,
     sub_550_2_n_20, sub_550_2_n_21, sub_550_2_n_22, sub_550_2_n_23,
     sub_550_2_n_24, sub_550_2_n_25, sub_550_2_n_26, sub_550_2_n_27,
     sub_550_2_n_28, sub_550_2_n_30, sub_550_2_n_38, sub_550_2_n_39,
     sub_550_2_n_40, sub_550_2_n_41, sub_550_2_n_43, sub_550_2_n_44,
     sub_550_2_n_45, sub_550_2_n_46, sub_550_2_n_48, sub_550_2_n_49,
     sub_550_2_n_50, sub_550_2_n_51, sub_550_2_n_52, sub_550_2_n_53,
     sub_550_2_n_54, sub_550_2_n_55, sub_550_2_n_56, sub_550_2_n_57,
     sub_550_2_n_58, sub_550_2_n_59, sub_550_2_n_60, sub_550_2_n_61,
     sub_550_2_n_62, sub_550_2_n_63, sub_550_2_n_64, sub_550_2_n_65,
     sub_550_2_n_66, sub_550_2_n_67, sub_550_2_n_68, sub_550_2_n_69,
     sub_550_2_n_70, sub_550_2_n_71, sub_550_2_n_72, sub_550_2_n_73,
     sub_550_2_n_74, sub_550_2_n_75, sub_550_2_n_76, sub_550_2_n_78,
     sub_550_2_n_79, sub_550_2_n_80, sub_550_2_n_81, sub_550_2_n_82,
     sub_550_2_n_83, sub_550_2_n_84, sub_550_2_n_85, sub_550_2_n_86,
     sub_550_2_n_87, sub_550_2_n_88, sub_550_2_n_89, sub_550_2_n_90,
     sub_550_2_n_91, sub_550_2_n_92, sub_550_2_n_93, sub_550_2_n_94,
     sub_550_2_n_95, sub_550_2_n_96, sub_550_2_n_97, sub_550_2_n_98,
     sub_550_2_n_99, sub_550_2_n_100, sub_550_2_n_101, sub_550_2_n_102,
     sub_550_2_n_103, sub_550_2_n_104, sub_550_2_n_105, sub_550_2_n_106,
     sub_550_2_n_107, sub_550_2_n_108, sub_550_2_n_109, sub_550_2_n_110,
     sub_550_2_n_111, sub_550_2_n_112, sub_550_2_n_113, sub_550_2_n_114,
     sub_550_2_n_115, sub_550_2_n_116, sub_550_2_n_117, sub_550_2_n_118,
     sub_550_2_n_119, sub_550_2_n_120, sub_550_2_n_122, sub_550_2_n_123,
     sub_550_2_n_124, sub_550_2_n_125, sub_550_2_n_126, sub_550_2_n_127,
     sub_550_2_n_128, sub_550_2_n_129, sub_550_2_n_130, sub_550_2_n_131,
     sub_550_2_n_132, sub_550_2_n_133, sub_550_2_n_134, sub_550_2_n_135,
     sub_550_2_n_136, sub_550_2_n_138, sub_550_2_n_139, sub_550_2_n_140,
     sub_550_2_n_141, sub_550_2_n_142, sub_550_2_n_144, sub_550_2_n_148,
     sub_571_2_n_0, sub_571_2_n_1, sub_571_2_n_2, sub_571_2_n_3, sub_571_2_n_4,
     sub_571_2_n_5, sub_571_2_n_6, sub_571_2_n_8, sub_571_2_n_9, sub_571_2_n_10,
     sub_571_2_n_11, sub_571_2_n_12, sub_571_2_n_13, sub_571_2_n_14,
     sub_571_2_n_15, sub_571_2_n_16, sub_571_2_n_17, sub_571_2_n_18,
     sub_571_2_n_19, sub_571_2_n_20, sub_571_2_n_21, sub_571_2_n_22,
     sub_571_2_n_23, sub_571_2_n_24, sub_571_2_n_25, sub_571_2_n_26,
     sub_571_2_n_27, sub_571_2_n_28, sub_571_2_n_29, sub_571_2_n_30,
     sub_571_2_n_38, sub_571_2_n_43, sub_571_2_n_44, sub_571_2_n_46,
     sub_571_2_n_47, sub_571_2_n_48, sub_571_2_n_51, sub_571_2_n_52,
     sub_571_2_n_54, sub_571_2_n_55, sub_571_2_n_56, sub_571_2_n_57,
     sub_571_2_n_58, sub_571_2_n_59, sub_571_2_n_60, sub_571_2_n_61,
     sub_571_2_n_62, sub_571_2_n_63, sub_571_2_n_64, sub_571_2_n_65,
     sub_571_2_n_66, sub_571_2_n_67, sub_571_2_n_68, sub_571_2_n_69,
     sub_571_2_n_70, sub_571_2_n_71, sub_571_2_n_72, sub_571_2_n_73,
     sub_571_2_n_74, sub_571_2_n_75, sub_571_2_n_76, sub_571_2_n_77,
     sub_571_2_n_78, sub_571_2_n_79, sub_571_2_n_80, sub_571_2_n_81,
     sub_571_2_n_82, sub_571_2_n_83, sub_571_2_n_84, sub_571_2_n_85,
     sub_571_2_n_86, sub_571_2_n_87, sub_571_2_n_89, sub_571_2_n_90,
     sub_571_2_n_91, sub_571_2_n_92, sub_571_2_n_93, sub_571_2_n_94,
     sub_571_2_n_95, sub_571_2_n_96, sub_571_2_n_97, sub_571_2_n_98,
     sub_571_2_n_99, sub_571_2_n_100, sub_571_2_n_101, sub_571_2_n_102,
     sub_571_2_n_103, sub_571_2_n_104, sub_571_2_n_105, sub_571_2_n_106,
     sub_571_2_n_107, sub_571_2_n_108, sub_571_2_n_109, sub_571_2_n_110,
     sub_571_2_n_111, sub_571_2_n_112, sub_571_2_n_113, sub_571_2_n_114,
     sub_571_2_n_115, sub_571_2_n_116, sub_571_2_n_117, sub_571_2_n_118,
     sub_571_2_n_119, sub_571_2_n_120, sub_571_2_n_121, sub_571_2_n_122,
     sub_571_2_n_123, sub_571_2_n_124, sub_571_2_n_125, sub_571_2_n_126,
     sub_571_2_n_127, sub_571_2_n_128, sub_571_2_n_129, sub_571_2_n_130,
     sub_571_2_n_131, sub_571_2_n_132, sub_571_2_n_133, sub_571_2_n_134,
     sub_571_2_n_135, sub_571_2_n_136, sub_571_2_n_137, sub_571_2_n_138,
     sub_571_2_n_139, sub_571_2_n_141, sub_571_2_n_142, sub_571_2_n_143,
     sub_571_2_n_146, sub_592_2_n_0, sub_592_2_n_1, sub_592_2_n_2, sub_592_2_n_3,
     sub_592_2_n_4, sub_592_2_n_5, sub_592_2_n_6, sub_592_2_n_7, sub_592_2_n_8,
     sub_592_2_n_9, sub_592_2_n_10, sub_592_2_n_11, sub_592_2_n_12,
     sub_592_2_n_13, sub_592_2_n_14, sub_592_2_n_15, sub_592_2_n_16,
     sub_592_2_n_17, sub_592_2_n_18, sub_592_2_n_19, sub_592_2_n_20,
     sub_592_2_n_21, sub_592_2_n_22, sub_592_2_n_23, sub_592_2_n_24,
     sub_592_2_n_25, sub_592_2_n_31, sub_592_2_n_36, sub_592_2_n_38,
     sub_592_2_n_43, sub_592_2_n_45, sub_592_2_n_46, sub_592_2_n_47,
     sub_592_2_n_48, sub_592_2_n_49, sub_592_2_n_50, sub_592_2_n_51,
     sub_592_2_n_53, sub_592_2_n_54, sub_592_2_n_55, sub_592_2_n_56,
     sub_592_2_n_57, sub_592_2_n_58, sub_592_2_n_59, sub_592_2_n_60,
     sub_592_2_n_61, sub_592_2_n_62, sub_592_2_n_63, sub_592_2_n_64,
     sub_592_2_n_65, sub_592_2_n_66, sub_592_2_n_67, sub_592_2_n_68,
     sub_592_2_n_69, sub_592_2_n_70, sub_592_2_n_71, sub_592_2_n_72,
     sub_592_2_n_73, sub_592_2_n_74, sub_592_2_n_75, sub_592_2_n_76,
     sub_592_2_n_77, sub_592_2_n_78, sub_592_2_n_79, sub_592_2_n_80,
     sub_592_2_n_81, sub_592_2_n_82, sub_592_2_n_83, sub_592_2_n_84,
     sub_592_2_n_85, sub_592_2_n_86, sub_592_2_n_87, sub_592_2_n_88,
     sub_592_2_n_89, sub_592_2_n_90, sub_592_2_n_91, sub_592_2_n_92,
     sub_592_2_n_94, sub_592_2_n_95, sub_592_2_n_96, sub_592_2_n_97,
     sub_592_2_n_98, sub_592_2_n_99, sub_592_2_n_100, sub_592_2_n_101,
     sub_592_2_n_102, sub_592_2_n_103, sub_592_2_n_104, sub_592_2_n_105,
     sub_592_2_n_106, sub_592_2_n_107, sub_592_2_n_108, sub_592_2_n_109,
     sub_592_2_n_110, sub_592_2_n_111, sub_592_2_n_112, sub_592_2_n_113,
     sub_592_2_n_114, sub_592_2_n_115, sub_592_2_n_116, sub_592_2_n_117,
     sub_592_2_n_118, sub_592_2_n_119, sub_592_2_n_120, sub_592_2_n_121,
     sub_592_2_n_122, sub_592_2_n_123, sub_592_2_n_124, sub_592_2_n_125,
     sub_592_2_n_126, sub_592_2_n_127, sub_592_2_n_128, sub_592_2_n_130,
     sub_592_2_n_131, sub_592_2_n_132, sub_592_2_n_133, sub_592_2_n_134,
     sub_592_2_n_135, sub_592_2_n_136, sub_592_2_n_137, sub_592_2_n_138,
     sub_592_2_n_139, sub_592_2_n_140, sub_592_2_n_141, sub_592_2_n_142,
     sub_592_2_n_143, sub_592_2_n_144, sub_592_2_n_145, sub_592_2_n_146,
     sub_592_2_n_147, sub_592_2_n_149, sub_592_2_n_150, sub_592_2_n_151,
     sub_592_2_n_152, sub_592_2_n_153, sub_592_2_n_154, sub_592_2_n_155,
     sub_592_2_n_156, sub_592_2_n_157, sub_592_2_n_158, sub_592_2_n_161,
     sub_592_2_n_162, sub_613_2_n_0, sub_613_2_n_1, sub_613_2_n_2, sub_613_2_n_3,
     sub_613_2_n_4, sub_613_2_n_5, sub_613_2_n_6, sub_613_2_n_7, sub_613_2_n_8,
     sub_613_2_n_9, sub_613_2_n_10, sub_613_2_n_12, sub_613_2_n_13,
     sub_613_2_n_14, sub_613_2_n_15, sub_613_2_n_16, sub_613_2_n_17,
     sub_613_2_n_18, sub_613_2_n_19, sub_613_2_n_20, sub_613_2_n_21,
     sub_613_2_n_22, sub_613_2_n_23, sub_613_2_n_24, sub_613_2_n_25,
     sub_613_2_n_31, sub_613_2_n_37, sub_613_2_n_40, sub_613_2_n_42,
     sub_613_2_n_43, sub_613_2_n_44, sub_613_2_n_45, sub_613_2_n_46,
     sub_613_2_n_47, sub_613_2_n_48, sub_613_2_n_50, sub_613_2_n_51,
     sub_613_2_n_52, sub_613_2_n_53, sub_613_2_n_54, sub_613_2_n_55,
     sub_613_2_n_56, sub_613_2_n_57, sub_613_2_n_58, sub_613_2_n_59,
     sub_613_2_n_60, sub_613_2_n_61, sub_613_2_n_62, sub_613_2_n_63,
     sub_613_2_n_64, sub_613_2_n_65, sub_613_2_n_66, sub_613_2_n_67,
     sub_613_2_n_68, sub_613_2_n_69, sub_613_2_n_70, sub_613_2_n_71,
     sub_613_2_n_72, sub_613_2_n_73, sub_613_2_n_74, sub_613_2_n_75,
     sub_613_2_n_76, sub_613_2_n_77, sub_613_2_n_78, sub_613_2_n_79,
     sub_613_2_n_80, sub_613_2_n_81, sub_613_2_n_82, sub_613_2_n_83,
     sub_613_2_n_84, sub_613_2_n_85, sub_613_2_n_86, sub_613_2_n_87,
     sub_613_2_n_88, sub_613_2_n_89, sub_613_2_n_90, sub_613_2_n_91,
     sub_613_2_n_92, sub_613_2_n_93, sub_613_2_n_95, sub_613_2_n_96,
     sub_613_2_n_97, sub_613_2_n_98, sub_613_2_n_99, sub_613_2_n_100,
     sub_613_2_n_101, sub_613_2_n_102, sub_613_2_n_103, sub_613_2_n_104,
     sub_613_2_n_105, sub_613_2_n_106, sub_613_2_n_107, sub_613_2_n_108,
     sub_613_2_n_109, sub_613_2_n_110, sub_613_2_n_111, sub_613_2_n_112,
     sub_613_2_n_113, sub_613_2_n_114, sub_613_2_n_115, sub_613_2_n_116,
     sub_613_2_n_117, sub_613_2_n_118, sub_613_2_n_119, sub_613_2_n_120,
     sub_613_2_n_121, sub_613_2_n_122, sub_613_2_n_123, sub_613_2_n_124,
     sub_613_2_n_125, sub_613_2_n_126, sub_613_2_n_127, sub_613_2_n_128,
     sub_613_2_n_129, sub_613_2_n_130, sub_613_2_n_131, sub_613_2_n_132,
     sub_613_2_n_133, sub_613_2_n_134, sub_613_2_n_135, sub_613_2_n_136,
     sub_613_2_n_137, sub_613_2_n_138, sub_613_2_n_139, sub_613_2_n_140,
     sub_613_2_n_141, sub_613_2_n_142, sub_613_2_n_143, sub_613_2_n_144,
     sub_613_2_n_145, sub_613_2_n_146, sub_613_2_n_147, sub_613_2_n_148,
     sub_613_2_n_149, sub_613_2_n_150, sub_613_2_n_151, sub_613_2_n_152,
     sub_613_2_n_153, sub_613_2_n_154, sub_613_2_n_155, sub_613_2_n_157,
     sub_613_2_n_158, sub_613_2_n_159, sub_613_2_n_160, sub_613_2_n_161,
     sub_613_2_n_162, sub_613_2_n_164, sub_613_2_n_165, sub_613_2_n_166,
     sub_613_2_n_167, sub_613_2_n_168, sub_613_2_n_169, sub_613_2_n_171,
     sub_613_2_n_172, sub_613_2_n_173, sub_613_2_n_176, sub_634_2_n_0,
     sub_634_2_n_1, sub_634_2_n_2, sub_634_2_n_3, sub_634_2_n_4, sub_634_2_n_5,
     sub_634_2_n_6, sub_634_2_n_7, sub_634_2_n_8, sub_634_2_n_9, sub_634_2_n_10,
     sub_634_2_n_11, sub_634_2_n_12, sub_634_2_n_13, sub_634_2_n_14,
     sub_634_2_n_15, sub_634_2_n_16, sub_634_2_n_17, sub_634_2_n_18,
     sub_634_2_n_19, sub_634_2_n_20, sub_634_2_n_21, sub_634_2_n_22,
     sub_634_2_n_23, sub_634_2_n_24, sub_634_2_n_25, sub_634_2_n_26,
     sub_634_2_n_27, sub_634_2_n_28, sub_634_2_n_32, sub_634_2_n_38,
     sub_634_2_n_40, sub_634_2_n_43, sub_634_2_n_44, sub_634_2_n_45,
     sub_634_2_n_46, sub_634_2_n_49, sub_634_2_n_50, sub_634_2_n_51,
     sub_634_2_n_52, sub_634_2_n_54, sub_634_2_n_55, sub_634_2_n_56,
     sub_634_2_n_57, sub_634_2_n_58, sub_634_2_n_59, sub_634_2_n_60,
     sub_634_2_n_61, sub_634_2_n_62, sub_634_2_n_63, sub_634_2_n_64,
     sub_634_2_n_65, sub_634_2_n_66, sub_634_2_n_67, sub_634_2_n_68,
     sub_634_2_n_69, sub_634_2_n_70, sub_634_2_n_71, sub_634_2_n_72,
     sub_634_2_n_73, sub_634_2_n_74, sub_634_2_n_75, sub_634_2_n_76,
     sub_634_2_n_77, sub_634_2_n_78, sub_634_2_n_79, sub_634_2_n_80,
     sub_634_2_n_81, sub_634_2_n_82, sub_634_2_n_83, sub_634_2_n_84,
     sub_634_2_n_85, sub_634_2_n_86, sub_634_2_n_87, sub_634_2_n_88,
     sub_634_2_n_89, sub_634_2_n_90, sub_634_2_n_91, sub_634_2_n_92,
     sub_634_2_n_93, sub_634_2_n_94, sub_634_2_n_95, sub_634_2_n_97,
     sub_634_2_n_98, sub_634_2_n_99, sub_634_2_n_100, sub_634_2_n_101,
     sub_634_2_n_102, sub_634_2_n_103, sub_634_2_n_104, sub_634_2_n_105,
     sub_634_2_n_106, sub_634_2_n_107, sub_634_2_n_108, sub_634_2_n_109,
     sub_634_2_n_110, sub_634_2_n_111, sub_634_2_n_112, sub_634_2_n_113,
     sub_634_2_n_114, sub_634_2_n_115, sub_634_2_n_116, sub_634_2_n_117,
     sub_634_2_n_118, sub_634_2_n_119, sub_634_2_n_120, sub_634_2_n_121,
     sub_634_2_n_122, sub_634_2_n_123, sub_634_2_n_124, sub_634_2_n_125,
     sub_634_2_n_126, sub_634_2_n_127, sub_634_2_n_128, sub_634_2_n_129,
     sub_634_2_n_130, sub_634_2_n_131, sub_634_2_n_132, sub_634_2_n_133,
     sub_634_2_n_135, sub_634_2_n_136, sub_634_2_n_137, sub_634_2_n_138,
     sub_634_2_n_139, sub_634_2_n_140, sub_634_2_n_141, sub_634_2_n_142,
     sub_634_2_n_143, sub_634_2_n_144, sub_634_2_n_145, sub_634_2_n_146,
     sub_634_2_n_147, sub_634_2_n_148, sub_634_2_n_149, sub_634_2_n_150,
     sub_634_2_n_151, sub_634_2_n_153, sub_634_2_n_154, sub_634_2_n_155,
     sub_634_2_n_156, sub_634_2_n_157, sub_634_2_n_159, sub_634_2_n_160,
     sub_634_2_n_161, sub_634_2_n_165, sub_634_2_n_167, sub_634_2_n_168,
     sub_655_2_n_1, sub_655_2_n_2, sub_655_2_n_3, sub_655_2_n_4, sub_655_2_n_5,
     sub_655_2_n_6, sub_655_2_n_7, sub_655_2_n_8, sub_655_2_n_9, sub_655_2_n_10,
     sub_655_2_n_11, sub_655_2_n_12, sub_655_2_n_13, sub_655_2_n_14,
     sub_655_2_n_15, sub_655_2_n_16, sub_655_2_n_17, sub_655_2_n_18,
     sub_655_2_n_19, sub_655_2_n_20, sub_655_2_n_21, sub_655_2_n_22,
     sub_655_2_n_23, sub_655_2_n_24, sub_655_2_n_25, sub_655_2_n_26,
     sub_655_2_n_27, sub_655_2_n_28, sub_655_2_n_29, sub_655_2_n_37,
     sub_655_2_n_41, sub_655_2_n_43, sub_655_2_n_44, sub_655_2_n_45,
     sub_655_2_n_46, sub_655_2_n_47, sub_655_2_n_49, sub_655_2_n_51,
     sub_655_2_n_52, sub_655_2_n_53, sub_655_2_n_54, sub_655_2_n_55,
     sub_655_2_n_56, sub_655_2_n_57, sub_655_2_n_58, sub_655_2_n_59,
     sub_655_2_n_60, sub_655_2_n_61, sub_655_2_n_62, sub_655_2_n_63,
     sub_655_2_n_64, sub_655_2_n_65, sub_655_2_n_66, sub_655_2_n_67,
     sub_655_2_n_68, sub_655_2_n_69, sub_655_2_n_70, sub_655_2_n_71,
     sub_655_2_n_72, sub_655_2_n_73, sub_655_2_n_74, sub_655_2_n_75,
     sub_655_2_n_76, sub_655_2_n_77, sub_655_2_n_78, sub_655_2_n_79,
     sub_655_2_n_80, sub_655_2_n_81, sub_655_2_n_82, sub_655_2_n_83,
     sub_655_2_n_84, sub_655_2_n_85, sub_655_2_n_86, sub_655_2_n_87,
     sub_655_2_n_88, sub_655_2_n_89, sub_655_2_n_90, sub_655_2_n_91,
     sub_655_2_n_92, sub_655_2_n_93, sub_655_2_n_94, sub_655_2_n_95,
     sub_655_2_n_96, sub_655_2_n_97, sub_655_2_n_99, sub_655_2_n_100,
     sub_655_2_n_101, sub_655_2_n_102, sub_655_2_n_103, sub_655_2_n_104,
     sub_655_2_n_105, sub_655_2_n_106, sub_655_2_n_107, sub_655_2_n_108,
     sub_655_2_n_109, sub_655_2_n_110, sub_655_2_n_111, sub_655_2_n_112,
     sub_655_2_n_113, sub_655_2_n_114, sub_655_2_n_115, sub_655_2_n_116,
     sub_655_2_n_117, sub_655_2_n_118, sub_655_2_n_119, sub_655_2_n_120,
     sub_655_2_n_121, sub_655_2_n_122, sub_655_2_n_123, sub_655_2_n_124,
     sub_655_2_n_125, sub_655_2_n_126, sub_655_2_n_127, sub_655_2_n_128,
     sub_655_2_n_129, sub_655_2_n_130, sub_655_2_n_131, sub_655_2_n_132,
     sub_655_2_n_133, sub_655_2_n_134, sub_655_2_n_135, sub_655_2_n_136,
     sub_655_2_n_137, sub_655_2_n_138, sub_655_2_n_139, sub_655_2_n_140,
     sub_655_2_n_141, sub_655_2_n_142, sub_655_2_n_143, sub_655_2_n_144,
     sub_655_2_n_145, sub_655_2_n_146, sub_655_2_n_147, sub_655_2_n_148,
     sub_655_2_n_149, sub_655_2_n_150, sub_655_2_n_151, sub_655_2_n_153,
     sub_655_2_n_154, sub_655_2_n_155, sub_655_2_n_156, sub_655_2_n_158,
     sub_655_2_n_159, sub_655_2_n_160, sub_655_2_n_161, sub_655_2_n_163,
     sub_655_2_n_164, sub_655_2_n_165, sub_655_2_n_166, sub_655_2_n_167,
     sub_655_2_n_168, sub_655_2_n_170, sub_655_2_n_171, sub_655_2_n_173,
     sub_655_2_n_176, sub_655_2_n_177, sub_655_2_n_178, sub_676_2_n_0,
     sub_676_2_n_1, sub_676_2_n_2, sub_676_2_n_3, sub_676_2_n_4, sub_676_2_n_5,
     sub_676_2_n_6, sub_676_2_n_7, sub_676_2_n_8, sub_676_2_n_9, sub_676_2_n_10,
     sub_676_2_n_11, sub_676_2_n_12, sub_676_2_n_13, sub_676_2_n_14,
     sub_676_2_n_15, sub_676_2_n_16, sub_676_2_n_17, sub_676_2_n_18,
     sub_676_2_n_19, sub_676_2_n_20, sub_676_2_n_21, sub_676_2_n_22,
     sub_676_2_n_23, sub_676_2_n_24, sub_676_2_n_25, sub_676_2_n_26,
     sub_676_2_n_27, sub_676_2_n_28, sub_676_2_n_29, sub_676_2_n_30,
     sub_676_2_n_31, sub_676_2_n_32, sub_676_2_n_33, sub_676_2_n_38,
     sub_676_2_n_49, sub_676_2_n_50, sub_676_2_n_51, sub_676_2_n_53,
     sub_676_2_n_55, sub_676_2_n_56, sub_676_2_n_57, sub_676_2_n_58,
     sub_676_2_n_59, sub_676_2_n_60, sub_676_2_n_61, sub_676_2_n_62,
     sub_676_2_n_63, sub_676_2_n_64, sub_676_2_n_65, sub_676_2_n_66,
     sub_676_2_n_67, sub_676_2_n_68, sub_676_2_n_69, sub_676_2_n_70,
     sub_676_2_n_71, sub_676_2_n_72, sub_676_2_n_73, sub_676_2_n_74,
     sub_676_2_n_75, sub_676_2_n_76, sub_676_2_n_77, sub_676_2_n_78,
     sub_676_2_n_79, sub_676_2_n_80, sub_676_2_n_81, sub_676_2_n_82,
     sub_676_2_n_83, sub_676_2_n_84, sub_676_2_n_85, sub_676_2_n_86,
     sub_676_2_n_87, sub_676_2_n_88, sub_676_2_n_89, sub_676_2_n_90,
     sub_676_2_n_91, sub_676_2_n_92, sub_676_2_n_93, sub_676_2_n_94,
     sub_676_2_n_95, sub_676_2_n_96, sub_676_2_n_97, sub_676_2_n_98,
     sub_676_2_n_99, sub_676_2_n_100, sub_676_2_n_101, sub_676_2_n_102,
     sub_676_2_n_103, sub_676_2_n_105, sub_676_2_n_106, sub_676_2_n_107,
     sub_676_2_n_108, sub_676_2_n_109, sub_676_2_n_110, sub_676_2_n_111,
     sub_676_2_n_112, sub_676_2_n_113, sub_676_2_n_114, sub_676_2_n_115,
     sub_676_2_n_116, sub_676_2_n_117, sub_676_2_n_118, sub_676_2_n_119,
     sub_676_2_n_120, sub_676_2_n_121, sub_676_2_n_122, sub_676_2_n_123,
     sub_676_2_n_124, sub_676_2_n_125, sub_676_2_n_126, sub_676_2_n_127,
     sub_676_2_n_128, sub_676_2_n_129, sub_676_2_n_130, sub_676_2_n_131,
     sub_676_2_n_132, sub_676_2_n_133, sub_676_2_n_134, sub_676_2_n_135,
     sub_676_2_n_136, sub_676_2_n_137, sub_676_2_n_138, sub_676_2_n_139,
     sub_676_2_n_140, sub_676_2_n_141, sub_676_2_n_142, sub_676_2_n_143,
     sub_676_2_n_144, sub_676_2_n_145, sub_676_2_n_146, sub_676_2_n_147,
     sub_676_2_n_148, sub_676_2_n_149, sub_676_2_n_150, sub_676_2_n_152,
     sub_676_2_n_153, sub_676_2_n_154, sub_676_2_n_155, sub_676_2_n_156,
     sub_676_2_n_157, sub_676_2_n_158, sub_676_2_n_159, sub_676_2_n_160,
     sub_676_2_n_161, sub_676_2_n_162, sub_676_2_n_163, sub_676_2_n_165,
     sub_676_2_n_166, sub_676_2_n_168, sub_676_2_n_169, sub_676_2_n_170,
     sub_676_2_n_171, sub_676_2_n_172, sub_676_2_n_173, sub_676_2_n_174,
     sub_676_2_n_175, sub_676_2_n_176, sub_676_2_n_177, sub_676_2_n_178,
     sub_676_2_n_181, sub_676_2_n_183, sub_676_2_n_184, sub_676_2_n_185,
     sub_676_2_n_188, sub_697_2_n_0, sub_697_2_n_1, sub_697_2_n_2, sub_697_2_n_3,
     sub_697_2_n_4, sub_697_2_n_5, sub_697_2_n_6, sub_697_2_n_7, sub_697_2_n_8,
     sub_697_2_n_9, sub_697_2_n_10, sub_697_2_n_11, sub_697_2_n_12,
     sub_697_2_n_13, sub_697_2_n_14, sub_697_2_n_15, sub_697_2_n_16,
     sub_697_2_n_17, sub_697_2_n_18, sub_697_2_n_19, sub_697_2_n_20,
     sub_697_2_n_21, sub_697_2_n_22, sub_697_2_n_25, sub_697_2_n_29,
     sub_697_2_n_32, sub_697_2_n_35, sub_697_2_n_36, sub_697_2_n_40,
     sub_697_2_n_41, sub_697_2_n_42, sub_697_2_n_43, sub_697_2_n_44,
     sub_697_2_n_45, sub_697_2_n_46, sub_697_2_n_48, sub_697_2_n_49,
     sub_697_2_n_50, sub_697_2_n_51, sub_697_2_n_52, sub_697_2_n_53,
     sub_697_2_n_54, sub_697_2_n_55, sub_697_2_n_56, sub_697_2_n_57,
     sub_697_2_n_58, sub_697_2_n_59, sub_697_2_n_60, sub_697_2_n_61,
     sub_697_2_n_62, sub_697_2_n_63, sub_697_2_n_64, sub_697_2_n_65,
     sub_697_2_n_66, sub_697_2_n_67, sub_697_2_n_68, sub_697_2_n_69,
     sub_697_2_n_70, sub_697_2_n_71, sub_697_2_n_72, sub_697_2_n_73,
     sub_697_2_n_74, sub_697_2_n_75, sub_697_2_n_76, sub_697_2_n_77,
     sub_697_2_n_78, sub_697_2_n_79, sub_697_2_n_80, sub_697_2_n_81,
     sub_697_2_n_82, sub_697_2_n_83, sub_697_2_n_84, sub_697_2_n_85,
     sub_697_2_n_86, sub_697_2_n_87, sub_697_2_n_88, sub_697_2_n_89,
     sub_697_2_n_90, sub_697_2_n_91, sub_697_2_n_92, sub_697_2_n_93,
     sub_697_2_n_94, sub_697_2_n_95, sub_697_2_n_96, sub_697_2_n_97,
     sub_697_2_n_98, sub_697_2_n_99, sub_697_2_n_100, sub_697_2_n_101,
     sub_697_2_n_102, sub_697_2_n_103, sub_697_2_n_104, sub_697_2_n_106,
     sub_697_2_n_107, sub_697_2_n_108, sub_697_2_n_109, sub_697_2_n_110,
     sub_697_2_n_111, sub_697_2_n_112, sub_697_2_n_113, sub_697_2_n_114,
     sub_697_2_n_115, sub_697_2_n_116, sub_697_2_n_117, sub_697_2_n_118,
     sub_697_2_n_119, sub_697_2_n_120, sub_697_2_n_121, sub_697_2_n_122,
     sub_697_2_n_123, sub_697_2_n_124, sub_697_2_n_125, sub_697_2_n_126,
     sub_697_2_n_127, sub_697_2_n_128, sub_697_2_n_129, sub_697_2_n_130,
     sub_697_2_n_131, sub_697_2_n_132, sub_697_2_n_133, sub_697_2_n_134,
     sub_697_2_n_135, sub_697_2_n_136, sub_697_2_n_137, sub_697_2_n_138,
     sub_697_2_n_139, sub_697_2_n_140, sub_697_2_n_141, sub_697_2_n_142,
     sub_697_2_n_143, sub_697_2_n_144, sub_697_2_n_145, sub_697_2_n_146,
     sub_697_2_n_147, sub_697_2_n_148, sub_697_2_n_149, sub_697_2_n_150,
     sub_697_2_n_151, sub_697_2_n_152, sub_697_2_n_153, sub_697_2_n_154,
     sub_697_2_n_155, sub_697_2_n_156, sub_697_2_n_158, sub_697_2_n_159,
     sub_697_2_n_160, sub_697_2_n_161, sub_697_2_n_162, sub_697_2_n_163,
     sub_697_2_n_164, sub_697_2_n_165, sub_697_2_n_166, sub_697_2_n_167,
     sub_697_2_n_168, sub_697_2_n_170, sub_697_2_n_171, sub_697_2_n_172,
     sub_697_2_n_173, sub_697_2_n_175, sub_697_2_n_176, sub_697_2_n_178,
     sub_697_2_n_179, sub_697_2_n_180, sub_697_2_n_181, sub_697_2_n_182,
     sub_697_2_n_183, sub_697_2_n_184, sub_697_2_n_185, sub_697_2_n_187,
     sub_697_2_n_188, sub_697_2_n_189, sub_697_2_n_191, sub_697_2_n_192,
     sub_697_2_n_193, sub_697_2_n_194, sub_697_2_n_195, sub_697_2_n_196,
     sub_697_2_n_200, sub_697_2_n_201, sub_697_2_n_202, sub_697_2_n_203,
     sub_697_2_n_206, sub_718_2_n_0, sub_718_2_n_1, sub_718_2_n_2, sub_718_2_n_3,
     sub_718_2_n_4, sub_718_2_n_5, sub_718_2_n_6, sub_718_2_n_7, sub_718_2_n_8,
     sub_718_2_n_9, sub_718_2_n_10, sub_718_2_n_11, sub_718_2_n_12,
     sub_718_2_n_13, sub_718_2_n_14, sub_718_2_n_15, sub_718_2_n_16,
     sub_718_2_n_17, sub_718_2_n_18, sub_718_2_n_19, sub_718_2_n_20,
     sub_718_2_n_21, sub_718_2_n_22, sub_718_2_n_23, sub_718_2_n_24,
     sub_718_2_n_25, sub_718_2_n_26, sub_718_2_n_33, sub_718_2_n_42,
     sub_718_2_n_43, sub_718_2_n_44, sub_718_2_n_46, sub_718_2_n_49,
     sub_718_2_n_50, sub_718_2_n_51, sub_718_2_n_52, sub_718_2_n_53,
     sub_718_2_n_54, sub_718_2_n_55, sub_718_2_n_56, sub_718_2_n_57,
     sub_718_2_n_58, sub_718_2_n_59, sub_718_2_n_60, sub_718_2_n_61,
     sub_718_2_n_62, sub_718_2_n_63, sub_718_2_n_64, sub_718_2_n_65,
     sub_718_2_n_66, sub_718_2_n_67, sub_718_2_n_68, sub_718_2_n_69,
     sub_718_2_n_70, sub_718_2_n_71, sub_718_2_n_72, sub_718_2_n_73,
     sub_718_2_n_74, sub_718_2_n_75, sub_718_2_n_76, sub_718_2_n_77,
     sub_718_2_n_78, sub_718_2_n_79, sub_718_2_n_80, sub_718_2_n_81,
     sub_718_2_n_82, sub_718_2_n_83, sub_718_2_n_84, sub_718_2_n_85,
     sub_718_2_n_86, sub_718_2_n_87, sub_718_2_n_88, sub_718_2_n_89,
     sub_718_2_n_90, sub_718_2_n_91, sub_718_2_n_92, sub_718_2_n_93,
     sub_718_2_n_94, sub_718_2_n_95, sub_718_2_n_96, sub_718_2_n_97,
     sub_718_2_n_98, sub_718_2_n_99, sub_718_2_n_100, sub_718_2_n_101,
     sub_718_2_n_102, sub_718_2_n_103, sub_718_2_n_104, sub_718_2_n_105,
     sub_718_2_n_106, sub_718_2_n_107, sub_718_2_n_109, sub_718_2_n_110,
     sub_718_2_n_111, sub_718_2_n_112, sub_718_2_n_113, sub_718_2_n_114,
     sub_718_2_n_115, sub_718_2_n_116, sub_718_2_n_117, sub_718_2_n_118,
     sub_718_2_n_119, sub_718_2_n_120, sub_718_2_n_121, sub_718_2_n_122,
     sub_718_2_n_123, sub_718_2_n_124, sub_718_2_n_125, sub_718_2_n_126,
     sub_718_2_n_127, sub_718_2_n_128, sub_718_2_n_129, sub_718_2_n_130,
     sub_718_2_n_131, sub_718_2_n_132, sub_718_2_n_133, sub_718_2_n_134,
     sub_718_2_n_135, sub_718_2_n_136, sub_718_2_n_137, sub_718_2_n_138,
     sub_718_2_n_139, sub_718_2_n_140, sub_718_2_n_141, sub_718_2_n_142,
     sub_718_2_n_143, sub_718_2_n_144, sub_718_2_n_145, sub_718_2_n_146,
     sub_718_2_n_147, sub_718_2_n_148, sub_718_2_n_149, sub_718_2_n_150,
     sub_718_2_n_151, sub_718_2_n_152, sub_718_2_n_153, sub_718_2_n_154,
     sub_718_2_n_155, sub_718_2_n_156, sub_718_2_n_157, sub_718_2_n_158,
     sub_718_2_n_159, sub_718_2_n_160, sub_718_2_n_161, sub_718_2_n_162,
     sub_718_2_n_163, sub_718_2_n_164, sub_718_2_n_165, sub_718_2_n_166,
     sub_718_2_n_167, sub_718_2_n_168, sub_718_2_n_169, sub_718_2_n_170,
     sub_718_2_n_171, sub_718_2_n_172, sub_718_2_n_173, sub_718_2_n_174,
     sub_718_2_n_175, sub_718_2_n_177, sub_718_2_n_178, sub_718_2_n_179,
     sub_718_2_n_180, sub_718_2_n_181, sub_718_2_n_182, sub_718_2_n_183,
     sub_718_2_n_184, sub_718_2_n_185, sub_718_2_n_186, sub_718_2_n_189,
     sub_718_2_n_190, sub_718_2_n_191, sub_718_2_n_192, sub_718_2_n_193,
     sub_718_2_n_197, sub_718_2_n_198, sub_718_2_n_199, sub_718_2_n_200,
     sub_718_2_n_202, sub_739_2_n_0, sub_739_2_n_1, sub_739_2_n_2, sub_739_2_n_3,
     sub_739_2_n_4, sub_739_2_n_5, sub_739_2_n_6, sub_739_2_n_7, sub_739_2_n_8,
     sub_739_2_n_9, sub_739_2_n_10, sub_739_2_n_11, sub_739_2_n_12,
     sub_739_2_n_13, sub_739_2_n_14, sub_739_2_n_15, sub_739_2_n_16,
     sub_739_2_n_17, sub_739_2_n_18, sub_739_2_n_19, sub_739_2_n_20,
     sub_739_2_n_21, sub_739_2_n_22, sub_739_2_n_23, sub_739_2_n_24,
     sub_739_2_n_25, sub_739_2_n_26, sub_739_2_n_27, sub_739_2_n_28,
     sub_739_2_n_29, sub_739_2_n_30, sub_739_2_n_31, sub_739_2_n_32,
     sub_739_2_n_33, sub_739_2_n_43, sub_739_2_n_49, sub_739_2_n_50,
     sub_739_2_n_51, sub_739_2_n_53, sub_739_2_n_54, sub_739_2_n_55,
     sub_739_2_n_56, sub_739_2_n_57, sub_739_2_n_58, sub_739_2_n_59,
     sub_739_2_n_60, sub_739_2_n_61, sub_739_2_n_62, sub_739_2_n_63,
     sub_739_2_n_64, sub_739_2_n_65, sub_739_2_n_66, sub_739_2_n_67,
     sub_739_2_n_68, sub_739_2_n_69, sub_739_2_n_70, sub_739_2_n_71,
     sub_739_2_n_72, sub_739_2_n_73, sub_739_2_n_74, sub_739_2_n_75,
     sub_739_2_n_76, sub_739_2_n_77, sub_739_2_n_78, sub_739_2_n_79,
     sub_739_2_n_80, sub_739_2_n_81, sub_739_2_n_82, sub_739_2_n_83,
     sub_739_2_n_84, sub_739_2_n_85, sub_739_2_n_86, sub_739_2_n_87,
     sub_739_2_n_88, sub_739_2_n_89, sub_739_2_n_90, sub_739_2_n_91,
     sub_739_2_n_92, sub_739_2_n_93, sub_739_2_n_94, sub_739_2_n_95,
     sub_739_2_n_97, sub_739_2_n_98, sub_739_2_n_99, sub_739_2_n_100,
     sub_739_2_n_101, sub_739_2_n_102, sub_739_2_n_103, sub_739_2_n_104,
     sub_739_2_n_105, sub_739_2_n_106, sub_739_2_n_107, sub_739_2_n_108,
     sub_739_2_n_109, sub_739_2_n_110, sub_739_2_n_111, sub_739_2_n_112,
     sub_739_2_n_113, sub_739_2_n_114, sub_739_2_n_115, sub_739_2_n_116,
     sub_739_2_n_117, sub_739_2_n_118, sub_739_2_n_119, sub_739_2_n_120,
     sub_739_2_n_121, sub_739_2_n_122, sub_739_2_n_123, sub_739_2_n_124,
     sub_739_2_n_125, sub_739_2_n_126, sub_739_2_n_127, sub_739_2_n_128,
     sub_739_2_n_129, sub_739_2_n_130, sub_739_2_n_131, sub_739_2_n_132,
     sub_739_2_n_133, sub_739_2_n_135, sub_739_2_n_136, sub_739_2_n_137,
     sub_739_2_n_138, sub_739_2_n_139, sub_739_2_n_140, sub_739_2_n_141,
     sub_739_2_n_142, sub_739_2_n_143, sub_739_2_n_144, sub_739_2_n_145,
     sub_739_2_n_146, sub_739_2_n_147, sub_739_2_n_148, sub_739_2_n_150,
     sub_739_2_n_151, sub_739_2_n_152, sub_739_2_n_155, sub_739_2_n_156,
     sub_739_2_n_157, sub_739_2_n_158, sub_739_2_n_159, sub_739_2_n_160,
     sub_739_2_n_161, sub_739_2_n_163, sub_739_2_n_164, sub_739_2_n_165,
     sub_739_2_n_166, sub_739_2_n_167, sub_739_2_n_168, sub_739_2_n_170,
     sub_739_2_n_171, sub_739_2_n_173, sub_739_2_n_176, sub_739_2_n_177,
     sub_739_2_n_178, sub_739_2_n_179, sub_739_2_n_180, sub_760_2_n_0,
     sub_760_2_n_1, sub_760_2_n_2, sub_760_2_n_3, sub_760_2_n_4, sub_760_2_n_5,
     sub_760_2_n_6, sub_760_2_n_7, sub_760_2_n_8, sub_760_2_n_9, sub_760_2_n_10,
     sub_760_2_n_11, sub_760_2_n_12, sub_760_2_n_13, sub_760_2_n_14,
     sub_760_2_n_15, sub_760_2_n_16, sub_760_2_n_17, sub_760_2_n_18,
     sub_760_2_n_19, sub_760_2_n_20, sub_760_2_n_21, sub_760_2_n_22,
     sub_760_2_n_23, sub_760_2_n_24, sub_760_2_n_25, sub_760_2_n_26,
     sub_760_2_n_27, sub_760_2_n_28, sub_760_2_n_29, sub_760_2_n_30,
     sub_760_2_n_31, sub_760_2_n_34, sub_760_2_n_45, sub_760_2_n_48,
     sub_760_2_n_51, sub_760_2_n_52, sub_760_2_n_55, sub_760_2_n_56,
     sub_760_2_n_57, sub_760_2_n_58, sub_760_2_n_59, sub_760_2_n_60,
     sub_760_2_n_61, sub_760_2_n_62, sub_760_2_n_63, sub_760_2_n_64,
     sub_760_2_n_65, sub_760_2_n_66, sub_760_2_n_67, sub_760_2_n_68,
     sub_760_2_n_69, sub_760_2_n_70, sub_760_2_n_71, sub_760_2_n_72,
     sub_760_2_n_73, sub_760_2_n_74, sub_760_2_n_75, sub_760_2_n_76,
     sub_760_2_n_77, sub_760_2_n_78, sub_760_2_n_79, sub_760_2_n_80,
     sub_760_2_n_81, sub_760_2_n_82, sub_760_2_n_83, sub_760_2_n_84,
     sub_760_2_n_85, sub_760_2_n_86, sub_760_2_n_87, sub_760_2_n_88,
     sub_760_2_n_89, sub_760_2_n_90, sub_760_2_n_91, sub_760_2_n_92,
     sub_760_2_n_93, sub_760_2_n_95, sub_760_2_n_96, sub_760_2_n_97,
     sub_760_2_n_98, sub_760_2_n_99, sub_760_2_n_100, sub_760_2_n_101,
     sub_760_2_n_102, sub_760_2_n_103, sub_760_2_n_104, sub_760_2_n_105,
     sub_760_2_n_106, sub_760_2_n_107, sub_760_2_n_108, sub_760_2_n_109,
     sub_760_2_n_110, sub_760_2_n_111, sub_760_2_n_112, sub_760_2_n_113,
     sub_760_2_n_114, sub_760_2_n_115, sub_760_2_n_116, sub_760_2_n_117,
     sub_760_2_n_118, sub_760_2_n_119, sub_760_2_n_120, sub_760_2_n_121,
     sub_760_2_n_122, sub_760_2_n_123, sub_760_2_n_124, sub_760_2_n_125,
     sub_760_2_n_126, sub_760_2_n_127, sub_760_2_n_128, sub_760_2_n_129,
     sub_760_2_n_130, sub_760_2_n_131, sub_760_2_n_132, sub_760_2_n_133,
     sub_760_2_n_134, sub_760_2_n_135, sub_760_2_n_136, sub_760_2_n_138,
     sub_760_2_n_139, sub_760_2_n_140, sub_760_2_n_142, sub_760_2_n_143,
     sub_760_2_n_144, sub_760_2_n_145, sub_760_2_n_146, sub_760_2_n_147,
     sub_760_2_n_148, sub_760_2_n_149, sub_760_2_n_150, sub_760_2_n_151,
     sub_760_2_n_152, sub_760_2_n_153, sub_760_2_n_154, sub_760_2_n_155,
     sub_760_2_n_156, sub_760_2_n_157, sub_760_2_n_158, sub_760_2_n_160,
     sub_760_2_n_161, sub_760_2_n_162, sub_760_2_n_163, sub_760_2_n_164,
     sub_760_2_n_165, sub_760_2_n_166, sub_760_2_n_169, sub_760_2_n_170,
     sub_760_2_n_171, sub_760_2_n_172, sub_760_2_n_174, sub_781_2_n_0,
     sub_781_2_n_1, sub_781_2_n_2, sub_781_2_n_3, sub_781_2_n_4, sub_781_2_n_5,
     sub_781_2_n_6, sub_781_2_n_7, sub_781_2_n_8, sub_781_2_n_9, sub_781_2_n_10,
     sub_781_2_n_11, sub_781_2_n_12, sub_781_2_n_13, sub_781_2_n_14,
     sub_781_2_n_15, sub_781_2_n_18, sub_781_2_n_21, sub_781_2_n_31,
     sub_781_2_n_35, sub_781_2_n_36, sub_781_2_n_37, sub_781_2_n_38,
     sub_781_2_n_39, sub_781_2_n_40, sub_781_2_n_41, sub_781_2_n_42,
     sub_781_2_n_43, sub_781_2_n_44, sub_781_2_n_45, sub_781_2_n_46,
     sub_781_2_n_47, sub_781_2_n_48, sub_781_2_n_49, sub_781_2_n_50,
     sub_781_2_n_51, sub_781_2_n_52, sub_781_2_n_53, sub_781_2_n_54,
     sub_781_2_n_55, sub_781_2_n_56, sub_781_2_n_57, sub_781_2_n_58,
     sub_781_2_n_59, sub_781_2_n_60, sub_781_2_n_61, sub_781_2_n_62,
     sub_781_2_n_63, sub_781_2_n_64, sub_781_2_n_65, sub_781_2_n_66,
     sub_781_2_n_67, sub_781_2_n_68, sub_781_2_n_69, sub_781_2_n_70,
     sub_781_2_n_71, sub_781_2_n_72, sub_781_2_n_73, sub_781_2_n_74,
     sub_781_2_n_75, sub_781_2_n_76, sub_781_2_n_77, sub_781_2_n_78,
     sub_781_2_n_79, sub_781_2_n_80, sub_781_2_n_81, sub_781_2_n_82,
     sub_781_2_n_83, sub_781_2_n_84, sub_781_2_n_85, sub_781_2_n_86,
     sub_781_2_n_87, sub_781_2_n_89, sub_781_2_n_90, sub_781_2_n_91,
     sub_781_2_n_92, sub_781_2_n_93, sub_781_2_n_94, sub_781_2_n_95,
     sub_781_2_n_96, sub_781_2_n_97, sub_781_2_n_98, sub_781_2_n_99,
     sub_781_2_n_100, sub_781_2_n_101, sub_781_2_n_102, sub_781_2_n_103,
     sub_781_2_n_104, sub_781_2_n_105, sub_781_2_n_106, sub_781_2_n_107,
     sub_781_2_n_108, sub_781_2_n_109, sub_781_2_n_110, sub_781_2_n_111,
     sub_781_2_n_112, sub_781_2_n_113, sub_781_2_n_114, sub_781_2_n_115,
     sub_781_2_n_116, sub_781_2_n_117, sub_781_2_n_118, sub_781_2_n_119,
     sub_781_2_n_120, sub_781_2_n_121, sub_781_2_n_122, sub_781_2_n_123,
     sub_781_2_n_124, sub_781_2_n_125, sub_781_2_n_126, sub_781_2_n_127,
     sub_781_2_n_128, sub_781_2_n_129, sub_781_2_n_130, sub_781_2_n_131,
     sub_781_2_n_132, sub_781_2_n_133, sub_781_2_n_134, sub_781_2_n_135,
     sub_781_2_n_136, sub_781_2_n_137, sub_781_2_n_139, sub_781_2_n_140,
     sub_781_2_n_141, sub_781_2_n_142, sub_781_2_n_143, sub_781_2_n_144,
     sub_781_2_n_145, sub_781_2_n_146, sub_781_2_n_147, sub_781_2_n_149,
     sub_781_2_n_150, sub_781_2_n_151, sub_781_2_n_152, sub_781_2_n_153,
     sub_781_2_n_154, sub_781_2_n_156, sub_781_2_n_157, sub_781_2_n_158,
     sub_781_2_n_159, sub_781_2_n_160, sub_781_2_n_161, sub_781_2_n_162,
     sub_781_2_n_164, sub_781_2_n_165, sub_781_2_n_166, sub_781_2_n_167,
     sub_781_2_n_168, sub_781_2_n_169, sub_781_2_n_174, sub_781_2_n_175,
     sub_781_2_n_176, sub_781_2_n_177, sub_781_2_n_178, sub_802_2_n_0,
     sub_802_2_n_1, sub_802_2_n_2, sub_802_2_n_3, sub_802_2_n_4, sub_802_2_n_5,
     sub_802_2_n_6, sub_802_2_n_7, sub_802_2_n_8, sub_802_2_n_14, sub_802_2_n_15,
     sub_802_2_n_16, sub_802_2_n_17, sub_802_2_n_19, sub_802_2_n_20,
     sub_802_2_n_21, sub_802_2_n_22, sub_802_2_n_23, sub_802_2_n_24,
     sub_802_2_n_25, sub_802_2_n_26, sub_802_2_n_27, sub_802_2_n_28,
     sub_802_2_n_29, sub_802_2_n_30, sub_802_2_n_31, sub_802_2_n_32,
     sub_802_2_n_33, sub_802_2_n_34, sub_802_2_n_35, sub_802_2_n_36,
     sub_802_2_n_37, sub_802_2_n_38, sub_802_2_n_39, sub_802_2_n_40,
     sub_802_2_n_41, sub_802_2_n_42, sub_802_2_n_43, sub_802_2_n_44,
     sub_802_2_n_45, sub_802_2_n_46, sub_802_2_n_47, sub_802_2_n_48,
     sub_802_2_n_49, sub_802_2_n_50, sub_802_2_n_51, sub_802_2_n_52,
     sub_802_2_n_53, sub_802_2_n_54, sub_802_2_n_55, sub_802_2_n_56,
     sub_802_2_n_57, sub_802_2_n_58, sub_802_2_n_59, sub_802_2_n_60,
     sub_802_2_n_61, sub_802_2_n_62, sub_802_2_n_63, sub_802_2_n_64,
     sub_802_2_n_65, sub_802_2_n_66, sub_802_2_n_67, sub_802_2_n_68,
     sub_802_2_n_69, sub_802_2_n_70, sub_802_2_n_71, sub_802_2_n_72,
     sub_802_2_n_73, sub_802_2_n_74, sub_802_2_n_75, sub_802_2_n_76,
     sub_802_2_n_77, sub_802_2_n_78, sub_802_2_n_79, sub_802_2_n_80,
     sub_802_2_n_81, sub_802_2_n_82, sub_802_2_n_83, sub_802_2_n_84,
     sub_802_2_n_85, sub_802_2_n_87, sub_802_2_n_88, sub_802_2_n_89,
     sub_802_2_n_90, sub_802_2_n_91, sub_802_2_n_92, sub_802_2_n_93,
     sub_802_2_n_94, sub_802_2_n_95, sub_802_2_n_96, sub_802_2_n_97,
     sub_802_2_n_98, sub_802_2_n_99, sub_802_2_n_100, sub_802_2_n_101,
     sub_802_2_n_102, sub_802_2_n_103, sub_802_2_n_104, sub_802_2_n_105,
     sub_802_2_n_106, sub_802_2_n_107, sub_802_2_n_108, sub_802_2_n_109,
     sub_802_2_n_110, sub_802_2_n_111, sub_802_2_n_112, sub_802_2_n_113,
     sub_802_2_n_114, sub_802_2_n_115, sub_802_2_n_116, sub_802_2_n_117,
     sub_802_2_n_118, sub_802_2_n_119, sub_802_2_n_120, sub_802_2_n_121,
     sub_802_2_n_122, sub_802_2_n_123, sub_802_2_n_124, sub_802_2_n_125,
     sub_802_2_n_126, sub_802_2_n_127, sub_802_2_n_129, sub_802_2_n_130,
     sub_802_2_n_131, sub_802_2_n_132, sub_802_2_n_133, sub_802_2_n_134,
     sub_802_2_n_135, sub_802_2_n_136, sub_802_2_n_137, sub_802_2_n_139,
     sub_802_2_n_140, sub_802_2_n_141, sub_802_2_n_142, sub_802_2_n_143,
     sub_802_2_n_144, sub_802_2_n_146, sub_802_2_n_147, sub_802_2_n_148,
     sub_802_2_n_149, sub_802_2_n_150, sub_802_2_n_151, sub_802_2_n_152,
     sub_802_2_n_153, sub_802_2_n_154, sub_802_2_n_155, sub_802_2_n_156,
     sub_802_2_n_161, sub_802_2_n_162, sub_802_2_n_163, sub_802_2_n_164,
     sub_802_2_n_165, sub_802_2_n_166, sub_802_2_n_173, sub_802_2_n_174,
     sub_802_2_n_175, sub_802_2_n_177, sub_802_2_n_178, sub_802_2_n_182,
     sub_823_2_n_0, sub_823_2_n_1, sub_823_2_n_2, sub_823_2_n_3, sub_823_2_n_4,
     sub_823_2_n_5, sub_823_2_n_6, sub_823_2_n_7, sub_823_2_n_8, sub_823_2_n_9,
     sub_823_2_n_10, sub_823_2_n_11, sub_823_2_n_12, sub_823_2_n_13,
     sub_823_2_n_14, sub_823_2_n_15, sub_823_2_n_20, sub_823_2_n_24,
     sub_823_2_n_25, sub_823_2_n_29, sub_823_2_n_31, sub_823_2_n_34,
     sub_823_2_n_35, sub_823_2_n_36, sub_823_2_n_37, sub_823_2_n_39,
     sub_823_2_n_40, sub_823_2_n_42, sub_823_2_n_43, sub_823_2_n_44,
     sub_823_2_n_45, sub_823_2_n_46, sub_823_2_n_47, sub_823_2_n_48,
     sub_823_2_n_49, sub_823_2_n_50, sub_823_2_n_51, sub_823_2_n_52,
     sub_823_2_n_53, sub_823_2_n_54, sub_823_2_n_55, sub_823_2_n_56,
     sub_823_2_n_57, sub_823_2_n_58, sub_823_2_n_59, sub_823_2_n_60,
     sub_823_2_n_61, sub_823_2_n_62, sub_823_2_n_63, sub_823_2_n_64,
     sub_823_2_n_65, sub_823_2_n_66, sub_823_2_n_67, sub_823_2_n_68,
     sub_823_2_n_69, sub_823_2_n_70, sub_823_2_n_71, sub_823_2_n_72,
     sub_823_2_n_73, sub_823_2_n_74, sub_823_2_n_75, sub_823_2_n_76,
     sub_823_2_n_77, sub_823_2_n_78, sub_823_2_n_79, sub_823_2_n_80,
     sub_823_2_n_81, sub_823_2_n_82, sub_823_2_n_83, sub_823_2_n_84,
     sub_823_2_n_85, sub_823_2_n_86, sub_823_2_n_87, sub_823_2_n_88,
     sub_823_2_n_89, sub_823_2_n_90, sub_823_2_n_91, sub_823_2_n_93,
     sub_823_2_n_94, sub_823_2_n_95, sub_823_2_n_96, sub_823_2_n_97,
     sub_823_2_n_98, sub_823_2_n_99, sub_823_2_n_100, sub_823_2_n_101,
     sub_823_2_n_102, sub_823_2_n_103, sub_823_2_n_104, sub_823_2_n_105,
     sub_823_2_n_106, sub_823_2_n_107, sub_823_2_n_108, sub_823_2_n_109,
     sub_823_2_n_110, sub_823_2_n_111, sub_823_2_n_112, sub_823_2_n_113,
     sub_823_2_n_114, sub_823_2_n_115, sub_823_2_n_116, sub_823_2_n_117,
     sub_823_2_n_118, sub_823_2_n_119, sub_823_2_n_120, sub_823_2_n_121,
     sub_823_2_n_122, sub_823_2_n_123, sub_823_2_n_124, sub_823_2_n_125,
     sub_823_2_n_126, sub_823_2_n_127, sub_823_2_n_128, sub_823_2_n_129,
     sub_823_2_n_130, sub_823_2_n_131, sub_823_2_n_133, sub_823_2_n_134,
     sub_823_2_n_135, sub_823_2_n_136, sub_823_2_n_137, sub_823_2_n_138,
     sub_823_2_n_139, sub_823_2_n_140, sub_823_2_n_141, sub_823_2_n_142,
     sub_823_2_n_145, sub_823_2_n_146, sub_823_2_n_147, sub_823_2_n_148,
     sub_823_2_n_149, sub_823_2_n_151, sub_823_2_n_153, sub_823_2_n_154,
     sub_823_2_n_155, sub_823_2_n_157, sub_823_2_n_158, sub_823_2_n_159,
     sub_823_2_n_160, sub_823_2_n_161, sub_823_2_n_163, sub_823_2_n_164,
     sub_823_2_n_165, sub_823_2_n_166, sub_823_2_n_168, sub_823_2_n_170,
     sub_823_2_n_171, sub_823_2_n_172, sub_823_2_n_173, sub_844_2_n_0,
     sub_844_2_n_1, sub_844_2_n_2, sub_844_2_n_3, sub_844_2_n_4, sub_844_2_n_5,
     sub_844_2_n_6, sub_844_2_n_7, sub_844_2_n_8, sub_844_2_n_9, sub_844_2_n_10,
     sub_844_2_n_11, sub_844_2_n_12, sub_844_2_n_13, sub_844_2_n_14,
     sub_844_2_n_15, sub_844_2_n_16, sub_844_2_n_17, sub_844_2_n_20,
     sub_844_2_n_24, sub_844_2_n_35, sub_844_2_n_36, sub_844_2_n_39,
     sub_844_2_n_40, sub_844_2_n_41, sub_844_2_n_42, sub_844_2_n_43,
     sub_844_2_n_44, sub_844_2_n_45, sub_844_2_n_46, sub_844_2_n_47,
     sub_844_2_n_48, sub_844_2_n_49, sub_844_2_n_50, sub_844_2_n_51,
     sub_844_2_n_52, sub_844_2_n_53, sub_844_2_n_54, sub_844_2_n_55,
     sub_844_2_n_56, sub_844_2_n_57, sub_844_2_n_58, sub_844_2_n_59,
     sub_844_2_n_60, sub_844_2_n_61, sub_844_2_n_62, sub_844_2_n_63,
     sub_844_2_n_64, sub_844_2_n_65, sub_844_2_n_66, sub_844_2_n_67,
     sub_844_2_n_68, sub_844_2_n_69, sub_844_2_n_70, sub_844_2_n_71,
     sub_844_2_n_72, sub_844_2_n_73, sub_844_2_n_74, sub_844_2_n_75,
     sub_844_2_n_76, sub_844_2_n_77, sub_844_2_n_78, sub_844_2_n_79,
     sub_844_2_n_80, sub_844_2_n_81, sub_844_2_n_82, sub_844_2_n_83,
     sub_844_2_n_84, sub_844_2_n_85, sub_844_2_n_86, sub_844_2_n_87,
     sub_844_2_n_88, sub_844_2_n_89, sub_844_2_n_91, sub_844_2_n_92,
     sub_844_2_n_93, sub_844_2_n_94, sub_844_2_n_95, sub_844_2_n_96,
     sub_844_2_n_97, sub_844_2_n_98, sub_844_2_n_99, sub_844_2_n_100,
     sub_844_2_n_101, sub_844_2_n_102, sub_844_2_n_103, sub_844_2_n_104,
     sub_844_2_n_105, sub_844_2_n_106, sub_844_2_n_107, sub_844_2_n_108,
     sub_844_2_n_109, sub_844_2_n_110, sub_844_2_n_111, sub_844_2_n_112,
     sub_844_2_n_113, sub_844_2_n_114, sub_844_2_n_115, sub_844_2_n_116,
     sub_844_2_n_117, sub_844_2_n_118, sub_844_2_n_119, sub_844_2_n_120,
     sub_844_2_n_121, sub_844_2_n_122, sub_844_2_n_123, sub_844_2_n_124,
     sub_844_2_n_125, sub_844_2_n_126, sub_844_2_n_127, sub_844_2_n_128,
     sub_844_2_n_129, sub_844_2_n_130, sub_844_2_n_131, sub_844_2_n_132,
     sub_844_2_n_133, sub_844_2_n_135, sub_844_2_n_136, sub_844_2_n_137,
     sub_844_2_n_138, sub_844_2_n_139, sub_844_2_n_140, sub_844_2_n_141,
     sub_844_2_n_142, sub_844_2_n_144, sub_844_2_n_145, sub_844_2_n_146,
     sub_844_2_n_147, sub_844_2_n_148, sub_844_2_n_149, sub_844_2_n_150,
     sub_844_2_n_151, sub_844_2_n_152, sub_844_2_n_153, sub_844_2_n_154,
     sub_844_2_n_156, sub_844_2_n_157, sub_844_2_n_158, sub_844_2_n_159,
     sub_844_2_n_160, sub_844_2_n_161, sub_844_2_n_162, sub_844_2_n_166,
     sub_844_2_n_167, sub_844_2_n_168, sub_844_2_n_169, sub_844_2_n_171,
     sub_865_2_n_0, sub_865_2_n_1, sub_865_2_n_2, sub_865_2_n_3, sub_865_2_n_4,
     sub_865_2_n_5, sub_865_2_n_6, sub_865_2_n_7, sub_865_2_n_8, sub_865_2_n_9,
     sub_865_2_n_10, sub_865_2_n_11, sub_865_2_n_12, sub_865_2_n_13,
     sub_865_2_n_14, sub_865_2_n_15, sub_865_2_n_16, sub_865_2_n_17,
     sub_865_2_n_18, sub_865_2_n_19, sub_865_2_n_20, sub_865_2_n_21,
     sub_865_2_n_22, sub_865_2_n_23, sub_865_2_n_24, sub_865_2_n_25,
     sub_865_2_n_27, sub_865_2_n_38, sub_865_2_n_39, sub_865_2_n_43,
     sub_865_2_n_44, sub_865_2_n_49, sub_865_2_n_50, sub_865_2_n_51,
     sub_865_2_n_52, sub_865_2_n_53, sub_865_2_n_54, sub_865_2_n_55,
     sub_865_2_n_56, sub_865_2_n_57, sub_865_2_n_58, sub_865_2_n_59,
     sub_865_2_n_60, sub_865_2_n_61, sub_865_2_n_62, sub_865_2_n_63,
     sub_865_2_n_64, sub_865_2_n_65, sub_865_2_n_66, sub_865_2_n_67,
     sub_865_2_n_68, sub_865_2_n_69, sub_865_2_n_70, sub_865_2_n_71,
     sub_865_2_n_72, sub_865_2_n_73, sub_865_2_n_74, sub_865_2_n_75,
     sub_865_2_n_76, sub_865_2_n_77, sub_865_2_n_78, sub_865_2_n_79,
     sub_865_2_n_80, sub_865_2_n_81, sub_865_2_n_82, sub_865_2_n_83,
     sub_865_2_n_84, sub_865_2_n_85, sub_865_2_n_86, sub_865_2_n_87,
     sub_865_2_n_88, sub_865_2_n_90, sub_865_2_n_91, sub_865_2_n_92,
     sub_865_2_n_93, sub_865_2_n_94, sub_865_2_n_95, sub_865_2_n_96,
     sub_865_2_n_97, sub_865_2_n_98, sub_865_2_n_99, sub_865_2_n_100,
     sub_865_2_n_101, sub_865_2_n_102, sub_865_2_n_103, sub_865_2_n_104,
     sub_865_2_n_105, sub_865_2_n_106, sub_865_2_n_107, sub_865_2_n_108,
     sub_865_2_n_109, sub_865_2_n_110, sub_865_2_n_111, sub_865_2_n_112,
     sub_865_2_n_113, sub_865_2_n_114, sub_865_2_n_115, sub_865_2_n_116,
     sub_865_2_n_117, sub_865_2_n_118, sub_865_2_n_119, sub_865_2_n_120,
     sub_865_2_n_121, sub_865_2_n_122, sub_865_2_n_123, sub_865_2_n_124,
     sub_865_2_n_125, sub_865_2_n_126, sub_865_2_n_127, sub_865_2_n_128,
     sub_865_2_n_129, sub_865_2_n_130, sub_865_2_n_132, sub_865_2_n_133,
     sub_865_2_n_134, sub_865_2_n_135, sub_865_2_n_136, sub_865_2_n_137,
     sub_865_2_n_138, sub_865_2_n_139, sub_865_2_n_140, sub_865_2_n_142,
     sub_865_2_n_143, sub_865_2_n_144, sub_865_2_n_145, sub_865_2_n_146,
     sub_865_2_n_147, sub_865_2_n_148, sub_865_2_n_149, sub_865_2_n_150,
     sub_865_2_n_151, sub_865_2_n_152, sub_865_2_n_153, sub_865_2_n_155,
     sub_865_2_n_156, sub_865_2_n_157, sub_865_2_n_158, sub_865_2_n_159,
     sub_865_2_n_160, sub_865_2_n_161, sub_865_2_n_162, sub_865_2_n_163,
     sub_865_2_n_165, sub_865_2_n_168, sub_886_2_n_0, sub_886_2_n_2,
     sub_886_2_n_3, sub_886_2_n_4, sub_886_2_n_5, sub_886_2_n_6, sub_886_2_n_7,
     sub_886_2_n_8, sub_886_2_n_9, sub_886_2_n_10, sub_886_2_n_11,
     sub_886_2_n_20, sub_886_2_n_21, sub_886_2_n_27, sub_886_2_n_30,
     sub_886_2_n_33, sub_886_2_n_36, sub_886_2_n_37, sub_886_2_n_38,
     sub_886_2_n_39, sub_886_2_n_40, sub_886_2_n_41, sub_886_2_n_42,
     sub_886_2_n_43, sub_886_2_n_44, sub_886_2_n_45, sub_886_2_n_46,
     sub_886_2_n_47, sub_886_2_n_48, sub_886_2_n_49, sub_886_2_n_50,
     sub_886_2_n_51, sub_886_2_n_52, sub_886_2_n_53, sub_886_2_n_54,
     sub_886_2_n_55, sub_886_2_n_56, sub_886_2_n_57, sub_886_2_n_58,
     sub_886_2_n_59, sub_886_2_n_60, sub_886_2_n_61, sub_886_2_n_62,
     sub_886_2_n_63, sub_886_2_n_64, sub_886_2_n_65, sub_886_2_n_66,
     sub_886_2_n_67, sub_886_2_n_68, sub_886_2_n_69, sub_886_2_n_70,
     sub_886_2_n_71, sub_886_2_n_72, sub_886_2_n_73, sub_886_2_n_74,
     sub_886_2_n_75, sub_886_2_n_76, sub_886_2_n_77, sub_886_2_n_78,
     sub_886_2_n_79, sub_886_2_n_80, sub_886_2_n_81, sub_886_2_n_82,
     sub_886_2_n_83, sub_886_2_n_84, sub_886_2_n_85, sub_886_2_n_86,
     sub_886_2_n_87, sub_886_2_n_88, sub_886_2_n_90, sub_886_2_n_91,
     sub_886_2_n_92, sub_886_2_n_93, sub_886_2_n_94, sub_886_2_n_95,
     sub_886_2_n_96, sub_886_2_n_97, sub_886_2_n_98, sub_886_2_n_99,
     sub_886_2_n_100, sub_886_2_n_101, sub_886_2_n_102, sub_886_2_n_103,
     sub_886_2_n_104, sub_886_2_n_105, sub_886_2_n_106, sub_886_2_n_107,
     sub_886_2_n_108, sub_886_2_n_109, sub_886_2_n_110, sub_886_2_n_111,
     sub_886_2_n_112, sub_886_2_n_113, sub_886_2_n_114, sub_886_2_n_115,
     sub_886_2_n_116, sub_886_2_n_117, sub_886_2_n_118, sub_886_2_n_119,
     sub_886_2_n_120, sub_886_2_n_121, sub_886_2_n_122, sub_886_2_n_123,
     sub_886_2_n_124, sub_886_2_n_125, sub_886_2_n_126, sub_886_2_n_127,
     sub_886_2_n_128, sub_886_2_n_129, sub_886_2_n_130, sub_886_2_n_131,
     sub_886_2_n_132, sub_886_2_n_133, sub_886_2_n_134, sub_886_2_n_135,
     sub_886_2_n_136, sub_886_2_n_137, sub_886_2_n_138, sub_886_2_n_139,
     sub_886_2_n_140, sub_886_2_n_141, sub_886_2_n_143, sub_886_2_n_144,
     sub_886_2_n_145, sub_886_2_n_146, sub_886_2_n_147, sub_886_2_n_148,
     sub_886_2_n_149, sub_886_2_n_150, sub_886_2_n_151, sub_886_2_n_152,
     sub_886_2_n_153, sub_886_2_n_154, sub_886_2_n_155, sub_886_2_n_156,
     sub_886_2_n_157, sub_886_2_n_159, sub_886_2_n_160, sub_886_2_n_161,
     sub_886_2_n_162, sub_886_2_n_163, sub_886_2_n_164, sub_886_2_n_167,
     sub_886_2_n_168, sub_886_2_n_169, sub_886_2_n_170, sub_886_2_n_171,
     sub_886_2_n_172, sub_886_2_n_173, sub_886_2_n_174, sub_886_2_n_175,
     sub_886_2_n_176, sub_886_2_n_177, sub_886_2_n_178, sub_907_2_n_0,
     sub_907_2_n_1, sub_907_2_n_2, sub_907_2_n_3, sub_907_2_n_4, sub_907_2_n_5,
     sub_907_2_n_6, sub_907_2_n_7, sub_907_2_n_8, sub_907_2_n_9, sub_907_2_n_10,
     sub_907_2_n_11, sub_907_2_n_12, sub_907_2_n_13, sub_907_2_n_14,
     sub_907_2_n_15, sub_907_2_n_16, sub_907_2_n_17, sub_907_2_n_20,
     sub_907_2_n_23, sub_907_2_n_29, sub_907_2_n_33, sub_907_2_n_34,
     sub_907_2_n_38, sub_907_2_n_39, sub_907_2_n_40, sub_907_2_n_41,
     sub_907_2_n_42, sub_907_2_n_43, sub_907_2_n_44, sub_907_2_n_45,
     sub_907_2_n_46, sub_907_2_n_47, sub_907_2_n_48, sub_907_2_n_49,
     sub_907_2_n_50, sub_907_2_n_51, sub_907_2_n_52, sub_907_2_n_53,
     sub_907_2_n_54, sub_907_2_n_55, sub_907_2_n_56, sub_907_2_n_57,
     sub_907_2_n_58, sub_907_2_n_59, sub_907_2_n_60, sub_907_2_n_61,
     sub_907_2_n_62, sub_907_2_n_63, sub_907_2_n_64, sub_907_2_n_65,
     sub_907_2_n_66, sub_907_2_n_67, sub_907_2_n_68, sub_907_2_n_69,
     sub_907_2_n_70, sub_907_2_n_71, sub_907_2_n_72, sub_907_2_n_73,
     sub_907_2_n_74, sub_907_2_n_75, sub_907_2_n_76, sub_907_2_n_77,
     sub_907_2_n_78, sub_907_2_n_79, sub_907_2_n_80, sub_907_2_n_81,
     sub_907_2_n_82, sub_907_2_n_83, sub_907_2_n_84, sub_907_2_n_85,
     sub_907_2_n_86, sub_907_2_n_88, sub_907_2_n_89, sub_907_2_n_90,
     sub_907_2_n_91, sub_907_2_n_92, sub_907_2_n_93, sub_907_2_n_94,
     sub_907_2_n_95, sub_907_2_n_96, sub_907_2_n_97, sub_907_2_n_98,
     sub_907_2_n_99, sub_907_2_n_100, sub_907_2_n_101, sub_907_2_n_102,
     sub_907_2_n_103, sub_907_2_n_104, sub_907_2_n_105, sub_907_2_n_106,
     sub_907_2_n_107, sub_907_2_n_108, sub_907_2_n_109, sub_907_2_n_110,
     sub_907_2_n_111, sub_907_2_n_112, sub_907_2_n_113, sub_907_2_n_114,
     sub_907_2_n_115, sub_907_2_n_116, sub_907_2_n_117, sub_907_2_n_118,
     sub_907_2_n_119, sub_907_2_n_120, sub_907_2_n_121, sub_907_2_n_122,
     sub_907_2_n_123, sub_907_2_n_124, sub_907_2_n_125, sub_907_2_n_126,
     sub_907_2_n_127, sub_907_2_n_128, sub_907_2_n_129, sub_907_2_n_130,
     sub_907_2_n_131, sub_907_2_n_132, sub_907_2_n_133, sub_907_2_n_134,
     sub_907_2_n_135, sub_907_2_n_137, sub_907_2_n_138, sub_907_2_n_139,
     sub_907_2_n_140, sub_907_2_n_141, sub_907_2_n_142, sub_907_2_n_143,
     sub_907_2_n_145, sub_907_2_n_147, sub_907_2_n_148, sub_907_2_n_150,
     sub_907_2_n_151, sub_907_2_n_153, sub_907_2_n_154, sub_907_2_n_155,
     sub_907_2_n_156, sub_907_2_n_159, sub_907_2_n_160, sub_907_2_n_161,
     sub_907_2_n_163, sub_907_2_n_164, sub_907_2_n_165, sub_907_2_n_166,
     sub_907_2_n_167, sub_907_2_n_169, sub_928_2_n_0, sub_928_2_n_1,
     sub_928_2_n_2, sub_928_2_n_3, sub_928_2_n_4, sub_928_2_n_5, sub_928_2_n_6,
     sub_928_2_n_7, sub_928_2_n_8, sub_928_2_n_9, sub_928_2_n_10, sub_928_2_n_11,
     sub_928_2_n_12, sub_928_2_n_13, sub_928_2_n_14, sub_928_2_n_15,
     sub_928_2_n_16, sub_928_2_n_17, sub_928_2_n_18, sub_928_2_n_19,
     sub_928_2_n_20, sub_928_2_n_21, sub_928_2_n_22, sub_928_2_n_28,
     sub_928_2_n_29, sub_928_2_n_40, sub_928_2_n_41, sub_928_2_n_42,
     sub_928_2_n_45, sub_928_2_n_46, sub_928_2_n_47, sub_928_2_n_48,
     sub_928_2_n_49, sub_928_2_n_50, sub_928_2_n_51, sub_928_2_n_52,
     sub_928_2_n_53, sub_928_2_n_54, sub_928_2_n_55, sub_928_2_n_56,
     sub_928_2_n_57, sub_928_2_n_58, sub_928_2_n_59, sub_928_2_n_60,
     sub_928_2_n_61, sub_928_2_n_62, sub_928_2_n_63, sub_928_2_n_64,
     sub_928_2_n_65, sub_928_2_n_66, sub_928_2_n_67, sub_928_2_n_68,
     sub_928_2_n_69, sub_928_2_n_70, sub_928_2_n_71, sub_928_2_n_72,
     sub_928_2_n_73, sub_928_2_n_74, sub_928_2_n_75, sub_928_2_n_76,
     sub_928_2_n_77, sub_928_2_n_78, sub_928_2_n_79, sub_928_2_n_80,
     sub_928_2_n_81, sub_928_2_n_82, sub_928_2_n_83, sub_928_2_n_84,
     sub_928_2_n_85, sub_928_2_n_86, sub_928_2_n_87, sub_928_2_n_88,
     sub_928_2_n_89, sub_928_2_n_90, sub_928_2_n_91, sub_928_2_n_92,
     sub_928_2_n_93, sub_928_2_n_95, sub_928_2_n_96, sub_928_2_n_97,
     sub_928_2_n_98, sub_928_2_n_99, sub_928_2_n_100, sub_928_2_n_101,
     sub_928_2_n_102, sub_928_2_n_103, sub_928_2_n_104, sub_928_2_n_105,
     sub_928_2_n_106, sub_928_2_n_107, sub_928_2_n_108, sub_928_2_n_109,
     sub_928_2_n_110, sub_928_2_n_111, sub_928_2_n_112, sub_928_2_n_113,
     sub_928_2_n_114, sub_928_2_n_115, sub_928_2_n_116, sub_928_2_n_117,
     sub_928_2_n_118, sub_928_2_n_119, sub_928_2_n_120, sub_928_2_n_121,
     sub_928_2_n_122, sub_928_2_n_123, sub_928_2_n_124, sub_928_2_n_125,
     sub_928_2_n_126, sub_928_2_n_127, sub_928_2_n_129, sub_928_2_n_130,
     sub_928_2_n_131, sub_928_2_n_132, sub_928_2_n_133, sub_928_2_n_134,
     sub_928_2_n_135, sub_928_2_n_136, sub_928_2_n_137, sub_928_2_n_138,
     sub_928_2_n_139, sub_928_2_n_141, sub_928_2_n_142, sub_928_2_n_143,
     sub_928_2_n_144, sub_928_2_n_146, sub_928_2_n_147, sub_928_2_n_148,
     sub_928_2_n_149, sub_928_2_n_150, sub_928_2_n_151, sub_928_2_n_152,
     sub_928_2_n_153, sub_928_2_n_154, sub_928_2_n_155, sub_928_2_n_157,
     sub_928_2_n_159, sub_928_2_n_160, sub_928_2_n_161, sub_928_2_n_162,
     sub_928_2_n_163, sub_928_2_n_164, sub_928_2_n_167, sub_928_2_n_168,
     sub_928_2_n_169, sub_928_2_n_170, sub_928_2_n_171, sub_949_2_n_0,
     sub_949_2_n_1, sub_949_2_n_2, sub_949_2_n_3, sub_949_2_n_4, sub_949_2_n_5,
     sub_949_2_n_6, sub_949_2_n_7, sub_949_2_n_8, sub_949_2_n_9, sub_949_2_n_10,
     sub_949_2_n_11, sub_949_2_n_12, sub_949_2_n_13, sub_949_2_n_14,
     sub_949_2_n_15, sub_949_2_n_16, sub_949_2_n_17, sub_949_2_n_18,
     sub_949_2_n_19, sub_949_2_n_22, sub_949_2_n_35, sub_949_2_n_36,
     sub_949_2_n_37, sub_949_2_n_38, sub_949_2_n_43, sub_949_2_n_44,
     sub_949_2_n_45, sub_949_2_n_46, sub_949_2_n_47, sub_949_2_n_48,
     sub_949_2_n_49, sub_949_2_n_50, sub_949_2_n_51, sub_949_2_n_52,
     sub_949_2_n_53, sub_949_2_n_54, sub_949_2_n_55, sub_949_2_n_56,
     sub_949_2_n_57, sub_949_2_n_58, sub_949_2_n_59, sub_949_2_n_60,
     sub_949_2_n_61, sub_949_2_n_62, sub_949_2_n_63, sub_949_2_n_64,
     sub_949_2_n_65, sub_949_2_n_66, sub_949_2_n_67, sub_949_2_n_68,
     sub_949_2_n_69, sub_949_2_n_70, sub_949_2_n_71, sub_949_2_n_72,
     sub_949_2_n_73, sub_949_2_n_74, sub_949_2_n_75, sub_949_2_n_76,
     sub_949_2_n_77, sub_949_2_n_78, sub_949_2_n_79, sub_949_2_n_80,
     sub_949_2_n_81, sub_949_2_n_82, sub_949_2_n_83, sub_949_2_n_84,
     sub_949_2_n_85, sub_949_2_n_86, sub_949_2_n_87, sub_949_2_n_88,
     sub_949_2_n_89, sub_949_2_n_91, sub_949_2_n_92, sub_949_2_n_93,
     sub_949_2_n_94, sub_949_2_n_95, sub_949_2_n_96, sub_949_2_n_97,
     sub_949_2_n_98, sub_949_2_n_99, sub_949_2_n_100, sub_949_2_n_101,
     sub_949_2_n_102, sub_949_2_n_103, sub_949_2_n_104, sub_949_2_n_105,
     sub_949_2_n_106, sub_949_2_n_107, sub_949_2_n_108, sub_949_2_n_109,
     sub_949_2_n_110, sub_949_2_n_111, sub_949_2_n_112, sub_949_2_n_113,
     sub_949_2_n_114, sub_949_2_n_115, sub_949_2_n_116, sub_949_2_n_117,
     sub_949_2_n_118, sub_949_2_n_119, sub_949_2_n_120, sub_949_2_n_121,
     sub_949_2_n_122, sub_949_2_n_123, sub_949_2_n_124, sub_949_2_n_125,
     sub_949_2_n_126, sub_949_2_n_127, sub_949_2_n_128, sub_949_2_n_129,
     sub_949_2_n_130, sub_949_2_n_132, sub_949_2_n_133, sub_949_2_n_134,
     sub_949_2_n_135, sub_949_2_n_136, sub_949_2_n_137, sub_949_2_n_138,
     sub_949_2_n_139, sub_949_2_n_140, sub_949_2_n_141, sub_949_2_n_142,
     sub_949_2_n_143, sub_949_2_n_144, sub_949_2_n_146, sub_949_2_n_147,
     sub_949_2_n_148, sub_949_2_n_149, sub_949_2_n_150, sub_949_2_n_151,
     sub_949_2_n_152, sub_949_2_n_154, sub_949_2_n_155, sub_949_2_n_156,
     sub_949_2_n_157, sub_949_2_n_159, sub_949_2_n_160, sub_949_2_n_161,
     sub_949_2_n_162, sub_949_2_n_163, sub_949_2_n_164, sub_949_2_n_165,
     sub_949_2_n_166, sub_949_2_n_168, sub_949_2_n_170, sub_970_2_n_0,
     sub_970_2_n_1, sub_970_2_n_2, sub_970_2_n_3, sub_970_2_n_4, sub_970_2_n_5,
     sub_970_2_n_6, sub_970_2_n_8, sub_970_2_n_12, sub_970_2_n_16,
     sub_970_2_n_19, sub_970_2_n_21, sub_970_2_n_22, sub_970_2_n_24,
     sub_970_2_n_25, sub_970_2_n_26, sub_970_2_n_27, sub_970_2_n_28,
     sub_970_2_n_29, sub_970_2_n_30, sub_970_2_n_31, sub_970_2_n_32,
     sub_970_2_n_33, sub_970_2_n_34, sub_970_2_n_35, sub_970_2_n_36,
     sub_970_2_n_37, sub_970_2_n_38, sub_970_2_n_39, sub_970_2_n_40,
     sub_970_2_n_41, sub_970_2_n_42, sub_970_2_n_43, sub_970_2_n_44,
     sub_970_2_n_45, sub_970_2_n_46, sub_970_2_n_47, sub_970_2_n_48,
     sub_970_2_n_49, sub_970_2_n_50, sub_970_2_n_51, sub_970_2_n_52,
     sub_970_2_n_53, sub_970_2_n_54, sub_970_2_n_55, sub_970_2_n_56,
     sub_970_2_n_57, sub_970_2_n_58, sub_970_2_n_59, sub_970_2_n_60,
     sub_970_2_n_61, sub_970_2_n_62, sub_970_2_n_63, sub_970_2_n_64,
     sub_970_2_n_65, sub_970_2_n_66, sub_970_2_n_67, sub_970_2_n_68,
     sub_970_2_n_69, sub_970_2_n_70, sub_970_2_n_71, sub_970_2_n_72,
     sub_970_2_n_73, sub_970_2_n_74, sub_970_2_n_75, sub_970_2_n_76,
     sub_970_2_n_77, sub_970_2_n_78, sub_970_2_n_79, sub_970_2_n_80,
     sub_970_2_n_81, sub_970_2_n_82, sub_970_2_n_83, sub_970_2_n_84,
     sub_970_2_n_85, sub_970_2_n_86, sub_970_2_n_88, sub_970_2_n_89,
     sub_970_2_n_90, sub_970_2_n_91, sub_970_2_n_92, sub_970_2_n_93,
     sub_970_2_n_94, sub_970_2_n_95, sub_970_2_n_96, sub_970_2_n_97,
     sub_970_2_n_98, sub_970_2_n_99, sub_970_2_n_100, sub_970_2_n_101,
     sub_970_2_n_102, sub_970_2_n_103, sub_970_2_n_104, sub_970_2_n_105,
     sub_970_2_n_106, sub_970_2_n_107, sub_970_2_n_108, sub_970_2_n_109,
     sub_970_2_n_110, sub_970_2_n_111, sub_970_2_n_112, sub_970_2_n_113,
     sub_970_2_n_114, sub_970_2_n_115, sub_970_2_n_116, sub_970_2_n_117,
     sub_970_2_n_118, sub_970_2_n_119, sub_970_2_n_120, sub_970_2_n_121,
     sub_970_2_n_122, sub_970_2_n_123, sub_970_2_n_124, sub_970_2_n_125,
     sub_970_2_n_126, sub_970_2_n_127, sub_970_2_n_128, sub_970_2_n_129,
     sub_970_2_n_130, sub_970_2_n_131, sub_970_2_n_132, sub_970_2_n_133,
     sub_970_2_n_134, sub_970_2_n_135, sub_970_2_n_136, sub_970_2_n_137,
     sub_970_2_n_138, sub_970_2_n_140, sub_970_2_n_141, sub_970_2_n_142,
     sub_970_2_n_143, sub_970_2_n_144, sub_970_2_n_145, sub_970_2_n_146,
     sub_970_2_n_147, sub_970_2_n_149, sub_970_2_n_150, sub_970_2_n_151,
     sub_970_2_n_152, sub_970_2_n_153, sub_970_2_n_154, sub_970_2_n_155,
     sub_970_2_n_157, sub_970_2_n_158, sub_970_2_n_159, sub_970_2_n_160,
     sub_970_2_n_161, sub_970_2_n_162, sub_970_2_n_167, sub_970_2_n_168,
     sub_970_2_n_169, sub_970_2_n_170, sub_970_2_n_171, sub_970_2_n_173,
     sub_970_2_n_177, sub_970_2_n_178, sub_970_2_n_179, sub_970_2_n_180,
     sub_970_2_n_183, sub_991_2_n_0, sub_991_2_n_1, sub_991_2_n_2, sub_991_2_n_3,
     sub_991_2_n_4, sub_991_2_n_5, sub_991_2_n_6, sub_991_2_n_7, sub_991_2_n_8,
     sub_991_2_n_9, sub_991_2_n_10, sub_991_2_n_11, sub_991_2_n_12,
     sub_991_2_n_13, sub_991_2_n_14, sub_991_2_n_15, sub_991_2_n_16,
     sub_991_2_n_17, sub_991_2_n_18, sub_991_2_n_19, sub_991_2_n_20,
     sub_991_2_n_21, sub_991_2_n_22, sub_991_2_n_25, sub_991_2_n_32,
     sub_991_2_n_43, sub_991_2_n_44, sub_991_2_n_47, sub_991_2_n_48,
     sub_991_2_n_49, sub_991_2_n_50, sub_991_2_n_51, sub_991_2_n_52,
     sub_991_2_n_53, sub_991_2_n_54, sub_991_2_n_55, sub_991_2_n_56,
     sub_991_2_n_57, sub_991_2_n_58, sub_991_2_n_59, sub_991_2_n_60,
     sub_991_2_n_61, sub_991_2_n_62, sub_991_2_n_63, sub_991_2_n_64,
     sub_991_2_n_65, sub_991_2_n_66, sub_991_2_n_67, sub_991_2_n_68,
     sub_991_2_n_69, sub_991_2_n_70, sub_991_2_n_71, sub_991_2_n_72,
     sub_991_2_n_73, sub_991_2_n_74, sub_991_2_n_75, sub_991_2_n_76,
     sub_991_2_n_77, sub_991_2_n_78, sub_991_2_n_79, sub_991_2_n_80,
     sub_991_2_n_81, sub_991_2_n_82, sub_991_2_n_83, sub_991_2_n_84,
     sub_991_2_n_85, sub_991_2_n_86, sub_991_2_n_87, sub_991_2_n_88,
     sub_991_2_n_89, sub_991_2_n_90, sub_991_2_n_91, sub_991_2_n_93,
     sub_991_2_n_94, sub_991_2_n_95, sub_991_2_n_96, sub_991_2_n_97,
     sub_991_2_n_98, sub_991_2_n_99, sub_991_2_n_100, sub_991_2_n_101,
     sub_991_2_n_102, sub_991_2_n_103, sub_991_2_n_104, sub_991_2_n_105,
     sub_991_2_n_106, sub_991_2_n_107, sub_991_2_n_108, sub_991_2_n_109,
     sub_991_2_n_110, sub_991_2_n_111, sub_991_2_n_112, sub_991_2_n_113,
     sub_991_2_n_114, sub_991_2_n_115, sub_991_2_n_116, sub_991_2_n_117,
     sub_991_2_n_118, sub_991_2_n_119, sub_991_2_n_120, sub_991_2_n_121,
     sub_991_2_n_122, sub_991_2_n_123, sub_991_2_n_124, sub_991_2_n_125,
     sub_991_2_n_126, sub_991_2_n_127, sub_991_2_n_128, sub_991_2_n_129,
     sub_991_2_n_130, sub_991_2_n_131, sub_991_2_n_132, sub_991_2_n_133,
     sub_991_2_n_135, sub_991_2_n_136, sub_991_2_n_137, sub_991_2_n_138,
     sub_991_2_n_139, sub_991_2_n_140, sub_991_2_n_141, sub_991_2_n_142,
     sub_991_2_n_143, sub_991_2_n_144, sub_991_2_n_145, sub_991_2_n_146,
     sub_991_2_n_147, sub_991_2_n_148, sub_991_2_n_150, sub_991_2_n_151,
     sub_991_2_n_152, sub_991_2_n_153, sub_991_2_n_154, sub_991_2_n_155,
     sub_991_2_n_156, sub_991_2_n_157, sub_991_2_n_158, sub_991_2_n_159,
     sub_991_2_n_161, sub_991_2_n_162, sub_991_2_n_163, sub_991_2_n_164,
     sub_991_2_n_165, sub_991_2_n_166, sub_991_2_n_167, sub_991_2_n_169,
     sub_991_2_n_170, sub_991_2_n_171, sub_991_2_n_172, sub_1012_2_n_0,
     sub_1012_2_n_2, sub_1012_2_n_3, sub_1012_2_n_4, sub_1012_2_n_5,
     sub_1012_2_n_6, sub_1012_2_n_7, sub_1012_2_n_8, sub_1012_2_n_9,
     sub_1012_2_n_23, sub_1012_2_n_24, sub_1012_2_n_25, sub_1012_2_n_27,
     sub_1012_2_n_28, sub_1012_2_n_29, sub_1012_2_n_30, sub_1012_2_n_31,
     sub_1012_2_n_32, sub_1012_2_n_33, sub_1012_2_n_34, sub_1012_2_n_35,
     sub_1012_2_n_36, sub_1012_2_n_37, sub_1012_2_n_38, sub_1012_2_n_39,
     sub_1012_2_n_40, sub_1012_2_n_41, sub_1012_2_n_42, sub_1012_2_n_43,
     sub_1012_2_n_44, sub_1012_2_n_45, sub_1012_2_n_46, sub_1012_2_n_47,
     sub_1012_2_n_48, sub_1012_2_n_49, sub_1012_2_n_50, sub_1012_2_n_51,
     sub_1012_2_n_52, sub_1012_2_n_53, sub_1012_2_n_54, sub_1012_2_n_55,
     sub_1012_2_n_56, sub_1012_2_n_57, sub_1012_2_n_58, sub_1012_2_n_59,
     sub_1012_2_n_60, sub_1012_2_n_61, sub_1012_2_n_62, sub_1012_2_n_63,
     sub_1012_2_n_64, sub_1012_2_n_65, sub_1012_2_n_66, sub_1012_2_n_67,
     sub_1012_2_n_68, sub_1012_2_n_69, sub_1012_2_n_70, sub_1012_2_n_71,
     sub_1012_2_n_72, sub_1012_2_n_73, sub_1012_2_n_74, sub_1012_2_n_75,
     sub_1012_2_n_76, sub_1012_2_n_77, sub_1012_2_n_78, sub_1012_2_n_79,
     sub_1012_2_n_80, sub_1012_2_n_81, sub_1012_2_n_82, sub_1012_2_n_83,
     sub_1012_2_n_84, sub_1012_2_n_85, sub_1012_2_n_86, sub_1012_2_n_87,
     sub_1012_2_n_88, sub_1012_2_n_89, sub_1012_2_n_90, sub_1012_2_n_91,
     sub_1012_2_n_93, sub_1012_2_n_94, sub_1012_2_n_95, sub_1012_2_n_96,
     sub_1012_2_n_97, sub_1012_2_n_98, sub_1012_2_n_99, sub_1012_2_n_100,
     sub_1012_2_n_101, sub_1012_2_n_102, sub_1012_2_n_103, sub_1012_2_n_104,
     sub_1012_2_n_105, sub_1012_2_n_106, sub_1012_2_n_107, sub_1012_2_n_108,
     sub_1012_2_n_109, sub_1012_2_n_110, sub_1012_2_n_111, sub_1012_2_n_112,
     sub_1012_2_n_113, sub_1012_2_n_114, sub_1012_2_n_115, sub_1012_2_n_116,
     sub_1012_2_n_117, sub_1012_2_n_118, sub_1012_2_n_119, sub_1012_2_n_120,
     sub_1012_2_n_121, sub_1012_2_n_122, sub_1012_2_n_123, sub_1012_2_n_124,
     sub_1012_2_n_125, sub_1012_2_n_126, sub_1012_2_n_127, sub_1012_2_n_128,
     sub_1012_2_n_129, sub_1012_2_n_130, sub_1012_2_n_131, sub_1012_2_n_132,
     sub_1012_2_n_133, sub_1012_2_n_134, sub_1012_2_n_135, sub_1012_2_n_136,
     sub_1012_2_n_137, sub_1012_2_n_138, sub_1012_2_n_140, sub_1012_2_n_141,
     sub_1012_2_n_142, sub_1012_2_n_143, sub_1012_2_n_144, sub_1012_2_n_145,
     sub_1012_2_n_147, sub_1012_2_n_148, sub_1012_2_n_149, sub_1012_2_n_151,
     sub_1012_2_n_152, sub_1012_2_n_153, sub_1012_2_n_154, sub_1012_2_n_155,
     sub_1012_2_n_156, sub_1012_2_n_157, sub_1012_2_n_159, sub_1012_2_n_160,
     sub_1012_2_n_161, sub_1012_2_n_162, sub_1012_2_n_163, sub_1012_2_n_164,
     sub_1012_2_n_165, sub_1012_2_n_166, sub_1012_2_n_167, sub_1012_2_n_168,
     sub_1012_2_n_169, sub_1012_2_n_170, sub_1012_2_n_174, sub_1012_2_n_175,
     sub_1012_2_n_176, sub_1012_2_n_177, sub_1012_2_n_178, sub_1012_2_n_179,
     sub_1012_2_n_180, sub_1012_2_n_181, sub_1012_2_n_184, sub_1012_2_n_185,
     sub_1012_2_n_186, sub_1012_2_n_187, sub_1012_2_n_188, sub_1033_2_n_0,
     sub_1033_2_n_1, sub_1033_2_n_2, sub_1033_2_n_3, sub_1033_2_n_4,
     sub_1033_2_n_5, sub_1033_2_n_6, sub_1033_2_n_7, sub_1033_2_n_8,
     sub_1033_2_n_9, sub_1033_2_n_10, sub_1033_2_n_11, sub_1033_2_n_12,
     sub_1033_2_n_13, sub_1033_2_n_16, sub_1033_2_n_22, sub_1033_2_n_29,
     sub_1033_2_n_31, sub_1033_2_n_32, sub_1033_2_n_34, sub_1033_2_n_35,
     sub_1033_2_n_36, sub_1033_2_n_37, sub_1033_2_n_38, sub_1033_2_n_39,
     sub_1033_2_n_40, sub_1033_2_n_41, sub_1033_2_n_42, sub_1033_2_n_43,
     sub_1033_2_n_44, sub_1033_2_n_45, sub_1033_2_n_46, sub_1033_2_n_47,
     sub_1033_2_n_48, sub_1033_2_n_49, sub_1033_2_n_50, sub_1033_2_n_51,
     sub_1033_2_n_52, sub_1033_2_n_53, sub_1033_2_n_54, sub_1033_2_n_55,
     sub_1033_2_n_56, sub_1033_2_n_57, sub_1033_2_n_58, sub_1033_2_n_59,
     sub_1033_2_n_60, sub_1033_2_n_61, sub_1033_2_n_62, sub_1033_2_n_63,
     sub_1033_2_n_64, sub_1033_2_n_65, sub_1033_2_n_66, sub_1033_2_n_67,
     sub_1033_2_n_68, sub_1033_2_n_69, sub_1033_2_n_70, sub_1033_2_n_71,
     sub_1033_2_n_72, sub_1033_2_n_73, sub_1033_2_n_74, sub_1033_2_n_75,
     sub_1033_2_n_76, sub_1033_2_n_77, sub_1033_2_n_78, sub_1033_2_n_79,
     sub_1033_2_n_81, sub_1033_2_n_82, sub_1033_2_n_83, sub_1033_2_n_84,
     sub_1033_2_n_85, sub_1033_2_n_86, sub_1033_2_n_87, sub_1033_2_n_88,
     sub_1033_2_n_89, sub_1033_2_n_90, sub_1033_2_n_91, sub_1033_2_n_92,
     sub_1033_2_n_93, sub_1033_2_n_94, sub_1033_2_n_95, sub_1033_2_n_96,
     sub_1033_2_n_97, sub_1033_2_n_98, sub_1033_2_n_99, sub_1033_2_n_100,
     sub_1033_2_n_101, sub_1033_2_n_102, sub_1033_2_n_103, sub_1033_2_n_104,
     sub_1033_2_n_105, sub_1033_2_n_106, sub_1033_2_n_107, sub_1033_2_n_108,
     sub_1033_2_n_109, sub_1033_2_n_110, sub_1033_2_n_111, sub_1033_2_n_112,
     sub_1033_2_n_113, sub_1033_2_n_114, sub_1033_2_n_115, sub_1033_2_n_116,
     sub_1033_2_n_117, sub_1033_2_n_118, sub_1033_2_n_119, sub_1033_2_n_120,
     sub_1033_2_n_121, sub_1033_2_n_123, sub_1033_2_n_124, sub_1033_2_n_125,
     sub_1033_2_n_126, sub_1033_2_n_127, sub_1033_2_n_128, sub_1033_2_n_129,
     sub_1033_2_n_130, sub_1033_2_n_132, sub_1033_2_n_133, sub_1033_2_n_134,
     sub_1033_2_n_135, sub_1033_2_n_136, sub_1033_2_n_137, sub_1033_2_n_138,
     sub_1033_2_n_139, sub_1033_2_n_140, sub_1033_2_n_142, sub_1033_2_n_143,
     sub_1033_2_n_145, sub_1033_2_n_146, sub_1033_2_n_147, sub_1033_2_n_148,
     sub_1033_2_n_149, sub_1033_2_n_151, sub_1033_2_n_152, sub_1033_2_n_153,
     sub_1033_2_n_154, sub_1033_2_n_156, sub_1033_2_n_157, sub_1033_2_n_158,
     sub_1033_2_n_160, sub_1033_2_n_163, sub_1033_2_n_164, sub_1033_2_n_165,
     sub_1033_2_n_166, sub_1033_2_n_167, sub_1054_2_n_0, sub_1054_2_n_1,
     sub_1054_2_n_2, sub_1054_2_n_3, sub_1054_2_n_4, sub_1054_2_n_5,
     sub_1054_2_n_6, sub_1054_2_n_7, sub_1054_2_n_8, sub_1054_2_n_10,
     sub_1054_2_n_20, sub_1054_2_n_21, sub_1054_2_n_23, sub_1054_2_n_24,
     sub_1054_2_n_28, sub_1054_2_n_29, sub_1054_2_n_30, sub_1054_2_n_31,
     sub_1054_2_n_32, sub_1054_2_n_33, sub_1054_2_n_34, sub_1054_2_n_35,
     sub_1054_2_n_36, sub_1054_2_n_37, sub_1054_2_n_38, sub_1054_2_n_39,
     sub_1054_2_n_40, sub_1054_2_n_41, sub_1054_2_n_42, sub_1054_2_n_43,
     sub_1054_2_n_44, sub_1054_2_n_45, sub_1054_2_n_46, sub_1054_2_n_47,
     sub_1054_2_n_48, sub_1054_2_n_49, sub_1054_2_n_50, sub_1054_2_n_51,
     sub_1054_2_n_52, sub_1054_2_n_53, sub_1054_2_n_54, sub_1054_2_n_55,
     sub_1054_2_n_56, sub_1054_2_n_57, sub_1054_2_n_58, sub_1054_2_n_59,
     sub_1054_2_n_60, sub_1054_2_n_61, sub_1054_2_n_62, sub_1054_2_n_63,
     sub_1054_2_n_64, sub_1054_2_n_65, sub_1054_2_n_66, sub_1054_2_n_67,
     sub_1054_2_n_68, sub_1054_2_n_69, sub_1054_2_n_70, sub_1054_2_n_71,
     sub_1054_2_n_72, sub_1054_2_n_74, sub_1054_2_n_75, sub_1054_2_n_76,
     sub_1054_2_n_77, sub_1054_2_n_78, sub_1054_2_n_79, sub_1054_2_n_80,
     sub_1054_2_n_81, sub_1054_2_n_82, sub_1054_2_n_83, sub_1054_2_n_84,
     sub_1054_2_n_85, sub_1054_2_n_86, sub_1054_2_n_87, sub_1054_2_n_88,
     sub_1054_2_n_89, sub_1054_2_n_90, sub_1054_2_n_91, sub_1054_2_n_92,
     sub_1054_2_n_93, sub_1054_2_n_94, sub_1054_2_n_95, sub_1054_2_n_96,
     sub_1054_2_n_97, sub_1054_2_n_98, sub_1054_2_n_99, sub_1054_2_n_100,
     sub_1054_2_n_101, sub_1054_2_n_102, sub_1054_2_n_103, sub_1054_2_n_104,
     sub_1054_2_n_105, sub_1054_2_n_106, sub_1054_2_n_107, sub_1054_2_n_108,
     sub_1054_2_n_109, sub_1054_2_n_110, sub_1054_2_n_111, sub_1054_2_n_112,
     sub_1054_2_n_113, sub_1054_2_n_114, sub_1054_2_n_115, sub_1054_2_n_116,
     sub_1054_2_n_117, sub_1054_2_n_118, sub_1054_2_n_119, sub_1054_2_n_120,
     sub_1054_2_n_121, sub_1054_2_n_122, sub_1054_2_n_123, sub_1054_2_n_124,
     sub_1054_2_n_125, sub_1054_2_n_126, sub_1054_2_n_127, sub_1054_2_n_129,
     sub_1054_2_n_130, sub_1054_2_n_131, sub_1054_2_n_132, sub_1054_2_n_133,
     sub_1054_2_n_134, sub_1054_2_n_136, sub_1054_2_n_137, sub_1054_2_n_139,
     sub_1054_2_n_140, sub_1054_2_n_141, sub_1054_2_n_143, sub_1054_2_n_144,
     sub_1054_2_n_146, sub_1054_2_n_147, sub_1054_2_n_148, sub_1054_2_n_149,
     sub_1054_2_n_151, sub_1054_2_n_152, sub_1054_2_n_154, sub_1054_2_n_155,
     sub_1054_2_n_156, sub_1054_2_n_157, sub_1054_2_n_158, sub_1054_2_n_159,
     sub_1054_2_n_162, sub_1054_2_n_163, sub_1054_2_n_164, sub_1054_2_n_166,
     sub_1054_2_n_167, sub_1075_2_n_0, sub_1075_2_n_1, sub_1075_2_n_2,
     sub_1075_2_n_3, sub_1075_2_n_4, sub_1075_2_n_5, sub_1075_2_n_6,
     sub_1075_2_n_7, sub_1075_2_n_8, sub_1075_2_n_17, sub_1075_2_n_20,
     sub_1075_2_n_22, sub_1075_2_n_23, sub_1075_2_n_24, sub_1075_2_n_25,
     sub_1075_2_n_26, sub_1075_2_n_27, sub_1075_2_n_28, sub_1075_2_n_29,
     sub_1075_2_n_30, sub_1075_2_n_31, sub_1075_2_n_32, sub_1075_2_n_33,
     sub_1075_2_n_34, sub_1075_2_n_35, sub_1075_2_n_36, sub_1075_2_n_37,
     sub_1075_2_n_38, sub_1075_2_n_39, sub_1075_2_n_40, sub_1075_2_n_41,
     sub_1075_2_n_42, sub_1075_2_n_43, sub_1075_2_n_44, sub_1075_2_n_45,
     sub_1075_2_n_46, sub_1075_2_n_47, sub_1075_2_n_48, sub_1075_2_n_49,
     sub_1075_2_n_50, sub_1075_2_n_51, sub_1075_2_n_52, sub_1075_2_n_53,
     sub_1075_2_n_54, sub_1075_2_n_55, sub_1075_2_n_56, sub_1075_2_n_57,
     sub_1075_2_n_58, sub_1075_2_n_59, sub_1075_2_n_60, sub_1075_2_n_61,
     sub_1075_2_n_62, sub_1075_2_n_63, sub_1075_2_n_64, sub_1075_2_n_65,
     sub_1075_2_n_66, sub_1075_2_n_67, sub_1075_2_n_68, sub_1075_2_n_69,
     sub_1075_2_n_70, sub_1075_2_n_71, sub_1075_2_n_72, sub_1075_2_n_73,
     sub_1075_2_n_74, sub_1075_2_n_75, sub_1075_2_n_76, sub_1075_2_n_77,
     sub_1075_2_n_78, sub_1075_2_n_79, sub_1075_2_n_81, sub_1075_2_n_82,
     sub_1075_2_n_83, sub_1075_2_n_84, sub_1075_2_n_85, sub_1075_2_n_86,
     sub_1075_2_n_87, sub_1075_2_n_88, sub_1075_2_n_89, sub_1075_2_n_90,
     sub_1075_2_n_91, sub_1075_2_n_92, sub_1075_2_n_93, sub_1075_2_n_94,
     sub_1075_2_n_95, sub_1075_2_n_96, sub_1075_2_n_97, sub_1075_2_n_98,
     sub_1075_2_n_99, sub_1075_2_n_100, sub_1075_2_n_101, sub_1075_2_n_102,
     sub_1075_2_n_103, sub_1075_2_n_104, sub_1075_2_n_105, sub_1075_2_n_106,
     sub_1075_2_n_107, sub_1075_2_n_108, sub_1075_2_n_109, sub_1075_2_n_110,
     sub_1075_2_n_111, sub_1075_2_n_112, sub_1075_2_n_113, sub_1075_2_n_114,
     sub_1075_2_n_115, sub_1075_2_n_116, sub_1075_2_n_117, sub_1075_2_n_118,
     sub_1075_2_n_119, sub_1075_2_n_120, sub_1075_2_n_121, sub_1075_2_n_122,
     sub_1075_2_n_123, sub_1075_2_n_124, sub_1075_2_n_125, sub_1075_2_n_126,
     sub_1075_2_n_127, sub_1075_2_n_128, sub_1075_2_n_129, sub_1075_2_n_130,
     sub_1075_2_n_131, sub_1075_2_n_132, sub_1075_2_n_133, sub_1075_2_n_135,
     sub_1075_2_n_136, sub_1075_2_n_137, sub_1075_2_n_138, sub_1075_2_n_139,
     sub_1075_2_n_140, sub_1075_2_n_141, sub_1075_2_n_143, sub_1075_2_n_144,
     sub_1075_2_n_145, sub_1075_2_n_148, sub_1075_2_n_149, sub_1075_2_n_152,
     sub_1075_2_n_153, sub_1075_2_n_154, sub_1075_2_n_156, sub_1075_2_n_157,
     sub_1075_2_n_158, sub_1075_2_n_159, sub_1075_2_n_160, sub_1075_2_n_161,
     sub_1075_2_n_162, sub_1075_2_n_163, sub_1075_2_n_164, sub_1075_2_n_165,
     sub_1075_2_n_167, sub_1075_2_n_168, sub_1075_2_n_169, sub_1075_2_n_170,
     sub_1075_2_n_171, sub_1075_2_n_172, sub_1075_2_n_173, sub_1075_2_n_177,
     sub_1075_2_n_178, sub_1075_2_n_179, sub_1075_2_n_181, sub_1075_2_n_182,
     sub_1075_2_n_183, sub_1096_2_n_0, sub_1096_2_n_1, sub_1096_2_n_2,
     sub_1096_2_n_3, sub_1096_2_n_4, sub_1096_2_n_6, sub_1096_2_n_8,
     sub_1096_2_n_9, sub_1096_2_n_10, sub_1096_2_n_11, sub_1096_2_n_12,
     sub_1096_2_n_13, sub_1096_2_n_14, sub_1096_2_n_15, sub_1096_2_n_16,
     sub_1096_2_n_17, sub_1096_2_n_18, sub_1096_2_n_19, sub_1096_2_n_20,
     sub_1096_2_n_21, sub_1096_2_n_22, sub_1096_2_n_23, sub_1096_2_n_24,
     sub_1096_2_n_25, sub_1096_2_n_26, sub_1096_2_n_27, sub_1096_2_n_28,
     sub_1096_2_n_29, sub_1096_2_n_30, sub_1096_2_n_31, sub_1096_2_n_32,
     sub_1096_2_n_33, sub_1096_2_n_34, sub_1096_2_n_35, sub_1096_2_n_36,
     sub_1096_2_n_37, sub_1096_2_n_38, sub_1096_2_n_39, sub_1096_2_n_40,
     sub_1096_2_n_41, sub_1096_2_n_42, sub_1096_2_n_43, sub_1096_2_n_44,
     sub_1096_2_n_45, sub_1096_2_n_46, sub_1096_2_n_47, sub_1096_2_n_48,
     sub_1096_2_n_49, sub_1096_2_n_50, sub_1096_2_n_51, sub_1096_2_n_52,
     sub_1096_2_n_53, sub_1096_2_n_54, sub_1096_2_n_55, sub_1096_2_n_56,
     sub_1096_2_n_57, sub_1096_2_n_58, sub_1096_2_n_59, sub_1096_2_n_60,
     sub_1096_2_n_61, sub_1096_2_n_62, sub_1096_2_n_63, sub_1096_2_n_64,
     sub_1096_2_n_65, sub_1096_2_n_67, sub_1096_2_n_68, sub_1096_2_n_69,
     sub_1096_2_n_70, sub_1096_2_n_71, sub_1096_2_n_72, sub_1096_2_n_73,
     sub_1096_2_n_74, sub_1096_2_n_75, sub_1096_2_n_76, sub_1096_2_n_77,
     sub_1096_2_n_78, sub_1096_2_n_79, sub_1096_2_n_80, sub_1096_2_n_81,
     sub_1096_2_n_82, sub_1096_2_n_83, sub_1096_2_n_84, sub_1096_2_n_85,
     sub_1096_2_n_86, sub_1096_2_n_87, sub_1096_2_n_88, sub_1096_2_n_89,
     sub_1096_2_n_90, sub_1096_2_n_91, sub_1096_2_n_92, sub_1096_2_n_93,
     sub_1096_2_n_94, sub_1096_2_n_95, sub_1096_2_n_96, sub_1096_2_n_97,
     sub_1096_2_n_98, sub_1096_2_n_99, sub_1096_2_n_100, sub_1096_2_n_101,
     sub_1096_2_n_102, sub_1096_2_n_103, sub_1096_2_n_104, sub_1096_2_n_105,
     sub_1096_2_n_106, sub_1096_2_n_107, sub_1096_2_n_108, sub_1096_2_n_109,
     sub_1096_2_n_110, sub_1096_2_n_111, sub_1096_2_n_113, sub_1096_2_n_114,
     sub_1096_2_n_115, sub_1096_2_n_116, sub_1096_2_n_118, sub_1096_2_n_119,
     sub_1096_2_n_120, sub_1096_2_n_121, sub_1096_2_n_124, sub_1096_2_n_125,
     sub_1096_2_n_126, sub_1096_2_n_127, sub_1096_2_n_128, sub_1096_2_n_131,
     sub_1096_2_n_132, sub_1096_2_n_134, sub_1096_2_n_135, sub_1096_2_n_136,
     sub_1096_2_n_137, sub_1096_2_n_138, sub_1096_2_n_140, sub_1096_2_n_141,
     sub_1096_2_n_142, sub_1096_2_n_143, sub_1096_2_n_144, sub_1096_2_n_149,
     sub_1096_2_n_150, sub_1096_2_n_151, sub_1096_2_n_152, sub_1096_2_n_153,
     sub_1096_2_n_154, sub_1096_2_n_155, sub_1096_2_n_163, sub_1096_2_n_164,
     sub_1096_2_n_165, sub_1096_2_n_166, sub_1096_2_n_169, sub_1117_2_n_0,
     sub_1117_2_n_1, sub_1117_2_n_2, sub_1117_2_n_3, sub_1117_2_n_4,
     sub_1117_2_n_5, sub_1117_2_n_6, sub_1117_2_n_7, sub_1117_2_n_8,
     sub_1117_2_n_9, sub_1117_2_n_10, sub_1117_2_n_11, sub_1117_2_n_12,
     sub_1117_2_n_13, sub_1117_2_n_14, sub_1117_2_n_15, sub_1117_2_n_16,
     sub_1117_2_n_17, sub_1117_2_n_18, sub_1117_2_n_19, sub_1117_2_n_20,
     sub_1117_2_n_21, sub_1117_2_n_22, sub_1117_2_n_23, sub_1117_2_n_24,
     sub_1117_2_n_25, sub_1117_2_n_26, sub_1117_2_n_27, sub_1117_2_n_28,
     sub_1117_2_n_29, sub_1117_2_n_30, sub_1117_2_n_31, sub_1117_2_n_32,
     sub_1117_2_n_33, sub_1117_2_n_34, sub_1117_2_n_35, sub_1117_2_n_36,
     sub_1117_2_n_37, sub_1117_2_n_38, sub_1117_2_n_39, sub_1117_2_n_40,
     sub_1117_2_n_41, sub_1117_2_n_42, sub_1117_2_n_43, sub_1117_2_n_44,
     sub_1117_2_n_45, sub_1117_2_n_46, sub_1117_2_n_47, sub_1117_2_n_48,
     sub_1117_2_n_49, sub_1117_2_n_50, sub_1117_2_n_51, sub_1117_2_n_52,
     sub_1117_2_n_53, sub_1117_2_n_54, sub_1117_2_n_55, sub_1117_2_n_56,
     sub_1117_2_n_57, sub_1117_2_n_58, sub_1117_2_n_59, sub_1117_2_n_60,
     sub_1117_2_n_61, sub_1117_2_n_62, sub_1117_2_n_64, sub_1117_2_n_65,
     sub_1117_2_n_66, sub_1117_2_n_67, sub_1117_2_n_68, sub_1117_2_n_69,
     sub_1117_2_n_70, sub_1117_2_n_71, sub_1117_2_n_72, sub_1117_2_n_73,
     sub_1117_2_n_74, sub_1117_2_n_75, sub_1117_2_n_76, sub_1117_2_n_77,
     sub_1117_2_n_78, sub_1117_2_n_79, sub_1117_2_n_80, sub_1117_2_n_81,
     sub_1117_2_n_82, sub_1117_2_n_83, sub_1117_2_n_84, sub_1117_2_n_85,
     sub_1117_2_n_86, sub_1117_2_n_87, sub_1117_2_n_88, sub_1117_2_n_89,
     sub_1117_2_n_90, sub_1117_2_n_91, sub_1117_2_n_92, sub_1117_2_n_93,
     sub_1117_2_n_94, sub_1117_2_n_95, sub_1117_2_n_96, sub_1117_2_n_97,
     sub_1117_2_n_98, sub_1117_2_n_99, sub_1117_2_n_100, sub_1117_2_n_101,
     sub_1117_2_n_102, sub_1117_2_n_103, sub_1117_2_n_104, sub_1117_2_n_105,
     sub_1117_2_n_107, sub_1117_2_n_108, sub_1117_2_n_109, sub_1117_2_n_111,
     sub_1117_2_n_112, sub_1117_2_n_113, sub_1117_2_n_114, sub_1117_2_n_117,
     sub_1117_2_n_118, sub_1117_2_n_119, sub_1117_2_n_122, sub_1117_2_n_124,
     sub_1117_2_n_125, sub_1117_2_n_126, sub_1117_2_n_127, sub_1117_2_n_129,
     sub_1117_2_n_133, sub_1117_2_n_134, sub_1117_2_n_135, sub_1117_2_n_136,
     sub_1117_2_n_137, sub_1117_2_n_139, sub_1117_2_n_140, sub_1117_2_n_141,
     sub_1117_2_n_146, sub_1117_2_n_150, sub_1117_2_n_151, sub_1117_2_n_152,
     sub_1117_2_n_157, sub_1138_2_n_0, sub_1138_2_n_1, sub_1138_2_n_2,
     sub_1138_2_n_3, sub_1138_2_n_4, sub_1138_2_n_5, sub_1138_2_n_6,
     sub_1138_2_n_7, sub_1138_2_n_8, sub_1138_2_n_9, sub_1138_2_n_10,
     sub_1138_2_n_11, sub_1138_2_n_12, sub_1138_2_n_13, sub_1138_2_n_14,
     sub_1138_2_n_15, sub_1138_2_n_16, sub_1138_2_n_17, sub_1138_2_n_18,
     sub_1138_2_n_19, sub_1138_2_n_20, sub_1138_2_n_21, sub_1138_2_n_22,
     sub_1138_2_n_23, sub_1138_2_n_24, sub_1138_2_n_25, sub_1138_2_n_26,
     sub_1138_2_n_27, sub_1138_2_n_28, sub_1138_2_n_29, sub_1138_2_n_30,
     sub_1138_2_n_31, sub_1138_2_n_32, sub_1138_2_n_33, sub_1138_2_n_34,
     sub_1138_2_n_35, sub_1138_2_n_36, sub_1138_2_n_37, sub_1138_2_n_38,
     sub_1138_2_n_39, sub_1138_2_n_40, sub_1138_2_n_41, sub_1138_2_n_42,
     sub_1138_2_n_43, sub_1138_2_n_44, sub_1138_2_n_45, sub_1138_2_n_46,
     sub_1138_2_n_47, sub_1138_2_n_48, sub_1138_2_n_49, sub_1138_2_n_50,
     sub_1138_2_n_51, sub_1138_2_n_52, sub_1138_2_n_53, sub_1138_2_n_54,
     sub_1138_2_n_55, sub_1138_2_n_56, sub_1138_2_n_57, sub_1138_2_n_58,
     sub_1138_2_n_59, sub_1138_2_n_60, sub_1138_2_n_62, sub_1138_2_n_63,
     sub_1138_2_n_64, sub_1138_2_n_65, sub_1138_2_n_66, sub_1138_2_n_67,
     sub_1138_2_n_68, sub_1138_2_n_69, sub_1138_2_n_70, sub_1138_2_n_71,
     sub_1138_2_n_72, sub_1138_2_n_73, sub_1138_2_n_74, sub_1138_2_n_75,
     sub_1138_2_n_76, sub_1138_2_n_77, sub_1138_2_n_78, sub_1138_2_n_79,
     sub_1138_2_n_80, sub_1138_2_n_81, sub_1138_2_n_82, sub_1138_2_n_83,
     sub_1138_2_n_84, sub_1138_2_n_85, sub_1138_2_n_86, sub_1138_2_n_87,
     sub_1138_2_n_88, sub_1138_2_n_89, sub_1138_2_n_90, sub_1138_2_n_91,
     sub_1138_2_n_92, sub_1138_2_n_93, sub_1138_2_n_94, sub_1138_2_n_95,
     sub_1138_2_n_96, sub_1138_2_n_97, sub_1138_2_n_98, sub_1138_2_n_99,
     sub_1138_2_n_100, sub_1138_2_n_102, sub_1138_2_n_103, sub_1138_2_n_104,
     sub_1138_2_n_105, sub_1138_2_n_107, sub_1138_2_n_108, sub_1138_2_n_111,
     sub_1138_2_n_112, sub_1138_2_n_113, sub_1138_2_n_114, sub_1138_2_n_117,
     sub_1138_2_n_118, sub_1138_2_n_120, sub_1138_2_n_121, sub_1138_2_n_122,
     sub_1138_2_n_123, sub_1138_2_n_125, sub_1138_2_n_130, sub_1138_2_n_131,
     sub_1138_2_n_132, sub_1138_2_n_133, sub_1138_2_n_134, sub_1138_2_n_135,
     sub_1138_2_n_143, sub_1138_2_n_144, sub_1138_2_n_145, sub_1138_2_n_146,
     sub_1138_2_n_151, sub_1159_2_n_0, sub_1159_2_n_1, sub_1159_2_n_2,
     sub_1159_2_n_3, sub_1159_2_n_4, sub_1159_2_n_5, sub_1159_2_n_6,
     sub_1159_2_n_7, sub_1159_2_n_8, sub_1159_2_n_9, sub_1159_2_n_10,
     sub_1159_2_n_11, sub_1159_2_n_12, sub_1159_2_n_13, sub_1159_2_n_14,
     sub_1159_2_n_15, sub_1159_2_n_16, sub_1159_2_n_17, sub_1159_2_n_18,
     sub_1159_2_n_19, sub_1159_2_n_20, sub_1159_2_n_21, sub_1159_2_n_22,
     sub_1159_2_n_23, sub_1159_2_n_24, sub_1159_2_n_25, sub_1159_2_n_26,
     sub_1159_2_n_27, sub_1159_2_n_28, sub_1159_2_n_29, sub_1159_2_n_30,
     sub_1159_2_n_31, sub_1159_2_n_32, sub_1159_2_n_33, sub_1159_2_n_34,
     sub_1159_2_n_35, sub_1159_2_n_36, sub_1159_2_n_37, sub_1159_2_n_38,
     sub_1159_2_n_39, sub_1159_2_n_40, sub_1159_2_n_41, sub_1159_2_n_42,
     sub_1159_2_n_43, sub_1159_2_n_44, sub_1159_2_n_45, sub_1159_2_n_46,
     sub_1159_2_n_47, sub_1159_2_n_48, sub_1159_2_n_49, sub_1159_2_n_50,
     sub_1159_2_n_51, sub_1159_2_n_52, sub_1159_2_n_53, sub_1159_2_n_54,
     sub_1159_2_n_55, sub_1159_2_n_56, sub_1159_2_n_57, sub_1159_2_n_58,
     sub_1159_2_n_59, sub_1159_2_n_61, sub_1159_2_n_62, sub_1159_2_n_63,
     sub_1159_2_n_64, sub_1159_2_n_65, sub_1159_2_n_66, sub_1159_2_n_67,
     sub_1159_2_n_68, sub_1159_2_n_69, sub_1159_2_n_70, sub_1159_2_n_71,
     sub_1159_2_n_72, sub_1159_2_n_73, sub_1159_2_n_74, sub_1159_2_n_75,
     sub_1159_2_n_76, sub_1159_2_n_77, sub_1159_2_n_78, sub_1159_2_n_79,
     sub_1159_2_n_80, sub_1159_2_n_81, sub_1159_2_n_82, sub_1159_2_n_83,
     sub_1159_2_n_84, sub_1159_2_n_85, sub_1159_2_n_86, sub_1159_2_n_87,
     sub_1159_2_n_88, sub_1159_2_n_89, sub_1159_2_n_90, sub_1159_2_n_91,
     sub_1159_2_n_92, sub_1159_2_n_93, sub_1159_2_n_94, sub_1159_2_n_95,
     sub_1159_2_n_96, sub_1159_2_n_98, sub_1159_2_n_99, sub_1159_2_n_100,
     sub_1159_2_n_101, sub_1159_2_n_103, sub_1159_2_n_104, sub_1159_2_n_107,
     sub_1159_2_n_108, sub_1159_2_n_109, sub_1159_2_n_112, sub_1159_2_n_113,
     sub_1159_2_n_115, sub_1159_2_n_116, sub_1159_2_n_117, sub_1159_2_n_118,
     sub_1159_2_n_120, sub_1159_2_n_124, sub_1159_2_n_125, sub_1159_2_n_126,
     sub_1159_2_n_127, sub_1159_2_n_129, sub_1159_2_n_130, sub_1159_2_n_131,
     sub_1159_2_n_136, sub_1159_2_n_140, sub_1159_2_n_141, sub_1159_2_n_142,
     sub_1159_2_n_147, sub_1180_2_n_0, sub_1180_2_n_1, sub_1180_2_n_2,
     sub_1180_2_n_3, sub_1180_2_n_4, sub_1180_2_n_5, sub_1180_2_n_6,
     sub_1180_2_n_7, sub_1180_2_n_8, sub_1180_2_n_9, sub_1180_2_n_10,
     sub_1180_2_n_11, sub_1180_2_n_12, sub_1180_2_n_13, sub_1180_2_n_14,
     sub_1180_2_n_15, sub_1180_2_n_16, sub_1180_2_n_17, sub_1180_2_n_18,
     sub_1180_2_n_19, sub_1180_2_n_20, sub_1180_2_n_21, sub_1180_2_n_22,
     sub_1180_2_n_23, sub_1180_2_n_24, sub_1180_2_n_25, sub_1180_2_n_26,
     sub_1180_2_n_27, sub_1180_2_n_28, sub_1180_2_n_29, sub_1180_2_n_30,
     sub_1180_2_n_31, sub_1180_2_n_32, sub_1180_2_n_33, sub_1180_2_n_34,
     sub_1180_2_n_35, sub_1180_2_n_36, sub_1180_2_n_37, sub_1180_2_n_38,
     sub_1180_2_n_39, sub_1180_2_n_40, sub_1180_2_n_41, sub_1180_2_n_42,
     sub_1180_2_n_43, sub_1180_2_n_44, sub_1180_2_n_45, sub_1180_2_n_46,
     sub_1180_2_n_47, sub_1180_2_n_48, sub_1180_2_n_49, sub_1180_2_n_50,
     sub_1180_2_n_51, sub_1180_2_n_52, sub_1180_2_n_53, sub_1180_2_n_54,
     sub_1180_2_n_55, sub_1180_2_n_56, sub_1180_2_n_57, sub_1180_2_n_58,
     sub_1180_2_n_59, sub_1180_2_n_61, sub_1180_2_n_62, sub_1180_2_n_63,
     sub_1180_2_n_64, sub_1180_2_n_65, sub_1180_2_n_66, sub_1180_2_n_67,
     sub_1180_2_n_68, sub_1180_2_n_69, sub_1180_2_n_70, sub_1180_2_n_71,
     sub_1180_2_n_72, sub_1180_2_n_73, sub_1180_2_n_74, sub_1180_2_n_75,
     sub_1180_2_n_76, sub_1180_2_n_77, sub_1180_2_n_78, sub_1180_2_n_79,
     sub_1180_2_n_80, sub_1180_2_n_81, sub_1180_2_n_82, sub_1180_2_n_83,
     sub_1180_2_n_84, sub_1180_2_n_85, sub_1180_2_n_86, sub_1180_2_n_87,
     sub_1180_2_n_88, sub_1180_2_n_89, sub_1180_2_n_90, sub_1180_2_n_91,
     sub_1180_2_n_92, sub_1180_2_n_93, sub_1180_2_n_94, sub_1180_2_n_95,
     sub_1180_2_n_96, sub_1180_2_n_97, sub_1180_2_n_99, sub_1180_2_n_100,
     sub_1180_2_n_101, sub_1180_2_n_102, sub_1180_2_n_104, sub_1180_2_n_105,
     sub_1180_2_n_108, sub_1180_2_n_109, sub_1180_2_n_110, sub_1180_2_n_113,
     sub_1180_2_n_114, sub_1180_2_n_116, sub_1180_2_n_117, sub_1180_2_n_118,
     sub_1180_2_n_119, sub_1180_2_n_121, sub_1180_2_n_125, sub_1180_2_n_126,
     sub_1180_2_n_127, sub_1180_2_n_128, sub_1180_2_n_130, sub_1180_2_n_131,
     sub_1180_2_n_132, sub_1180_2_n_137, sub_1180_2_n_141, sub_1180_2_n_142,
     sub_1180_2_n_143, sub_1180_2_n_148, sub_1199_2_n_0, sub_1199_2_n_1,
     sub_1199_2_n_3, sub_1199_2_n_4, sub_1199_2_n_5, sub_1199_2_n_6,
     sub_1199_2_n_7, sub_1199_2_n_8, sub_1199_2_n_9, sub_1199_2_n_10,
     sub_1199_2_n_11, sub_1199_2_n_12, sub_1199_2_n_13, sub_1199_2_n_14,
     sub_1199_2_n_15, sub_1199_2_n_16, sub_1199_2_n_17, sub_1199_2_n_18,
     sub_1199_2_n_19, sub_1199_2_n_20, sub_1199_2_n_21, sub_1199_2_n_22,
     sub_1199_2_n_23, sub_1199_2_n_24, sub_1199_2_n_25, sub_1199_2_n_26,
     sub_1199_2_n_27, sub_1199_2_n_28, sub_1199_2_n_29, sub_1199_2_n_30,
     sub_1199_2_n_31, sub_1199_2_n_32, sub_1199_2_n_33, sub_1199_2_n_34,
     sub_1199_2_n_35, sub_1199_2_n_36, sub_1199_2_n_37, sub_1199_2_n_38,
     sub_1199_2_n_39, sub_1199_2_n_40, sub_1199_2_n_41, sub_1199_2_n_42,
     sub_1199_2_n_43, sub_1199_2_n_44, sub_1199_2_n_45, sub_1199_2_n_46,
     sub_1199_2_n_47, sub_1199_2_n_48, sub_1199_2_n_49, sub_1199_2_n_50,
     sub_1199_2_n_51, sub_1199_2_n_52, sub_1199_2_n_53, sub_1199_2_n_54,
     sub_1199_2_n_55, sub_1199_2_n_56, sub_1199_2_n_57, sub_1199_2_n_58,
     sub_1199_2_n_59, sub_1199_2_n_60, sub_1199_2_n_61, sub_1199_2_n_62,
     sub_1199_2_n_63, sub_1199_2_n_64, sub_1199_2_n_65, sub_1199_2_n_66,
     sub_1199_2_n_67, sub_1199_2_n_68, sub_1199_2_n_69, sub_1199_2_n_70,
     sub_1199_2_n_71, sub_1199_2_n_72, sub_1199_2_n_73, sub_1199_2_n_74,
     sub_1199_2_n_75, sub_1199_2_n_76, sub_1199_2_n_77, sub_1199_2_n_78, stall,
     clk, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293,
     n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302,
     n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311,
     n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320,
     n_1321, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404,
     n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413,
     n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422,
     n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431,
     n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440,
     n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449,
     n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458,
     n_1459, n_1461, n_1462, n_1466, n_1467, n_1468, n_1470, n_1471, n_1472,
     n_1473, n_1474, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482,
     n_1484, n_1485, n_1486, n_1487, n_1488, n_1490, n_1491, n_1492, n_1493,
     n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502,
     n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1513,
     n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522,
     n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531,
     n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540,
     n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549,
     n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558,
     n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567,
     n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576,
     n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585,
     n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594,
     n_1595, n_1596, n_1597, n_1598, n_1599, asc001_0_0_, asc001_0_1_,
     asc001_0_2_, asc001_0_3_, asc001_0_4_, asc001_0_5_, asc001_0_6_,
     asc001_0_7_, asc001_0_8_, asc001_0_9_, asc001_0_10_, asc001_0_11_,
     asc001_0_12_, asc001_0_13_, asc001_0_14_, asc001_0_15_, asc001_0_16_,
     asc001_0_17_, asc001_0_18_, asc001_0_19_, asc001_0_20_, asc001_0_21_,
     asc001_0_22_, asc001_0_23_, asc001_0_24_, asc001_0_25_, asc001_0_26_,
     asc001_0_27_, asc001_0_28_, asc001_0_29_, asc001_0_30_, asc001_0_31_,
     asc001_0_32_, asc001_0_33_, asc001_0_34_, asc001_0_35_, asc001_0_36_,
     in1_1_0_, in1_1_24_, in1_2_0_, in1_4_0_, in1_4_1_, in1_4_24_, in1_5_0_,
     in1_5_1_, in1_7_0_, in1_7_1_, in1_7_2_, in1_7_24_, in1_8_0_, in1_8_1_,
     in1_8_2_, in1_10_0_, in1_10_1_, in1_10_2_, in1_10_3_, in1_10_24_, in1_11_0_,
     in1_11_1_, in1_11_2_, in1_11_3_, in1_13_0_, in1_13_1_, in1_13_2_, in1_13_3_,
     in1_13_4_, in1_13_24_, in1_14_0_, in1_14_1_, in1_14_2_, in1_14_3_,
     in1_14_4_, in1_16_0_, in1_16_1_, in1_16_2_, in1_16_3_, in1_16_4_, in1_16_5_,
     in1_16_24_, in1_17_0_, in1_17_1_, in1_17_2_, in1_17_3_, in1_17_4_,
     in1_17_5_, in1_19_0_, in1_19_1_, in1_19_2_, in1_19_3_, in1_19_4_, in1_19_5_,
     in1_19_6_, in1_19_24_, in1_20_0_, in1_20_1_, in1_20_2_, in1_20_3_,
     in1_20_4_, in1_20_5_, in1_20_6_, in1_22_0_, in1_22_1_, in1_22_2_, in1_22_3_,
     in1_22_4_, in1_22_5_, in1_22_6_, in1_22_7_, in1_22_24_, in1_23_0_,
     in1_23_1_, in1_23_2_, in1_23_3_, in1_23_4_, in1_23_5_, in1_23_6_, in1_23_7_,
     in1_25_0_, in1_25_1_, in1_25_2_, in1_25_3_, in1_25_4_, in1_25_5_, in1_25_6_,
     in1_25_7_, in1_25_8_, in1_25_24_, in1_26_0_, in1_26_1_, in1_26_2_,
     in1_26_3_, in1_26_4_, in1_26_5_, in1_26_6_, in1_26_7_, in1_26_8_, in1_28_0_,
     in1_28_1_, in1_28_2_, in1_28_3_, in1_28_4_, in1_28_5_, in1_28_6_, in1_28_7_,
     in1_28_8_, in1_28_9_, in1_28_24_, in1_29_0_, in1_29_1_, in1_29_2_,
     in1_29_3_, in1_29_4_, in1_29_5_, in1_29_6_, in1_29_7_, in1_29_8_, in1_29_9_,
     in1_31_0_, in1_31_1_, in1_31_2_, in1_31_3_, in1_31_4_, in1_31_5_, in1_31_6_,
     in1_31_7_, in1_31_8_, in1_31_9_, in1_31_10_, in1_31_24_, in1_32_0_,
     in1_32_1_, in1_32_2_, in1_32_3_, in1_32_4_, in1_32_5_, in1_32_6_, in1_32_7_,
     in1_32_8_, in1_32_9_, in1_32_10_, in1_34_0_, in1_34_1_, in1_34_2_,
     in1_34_3_, in1_34_4_, in1_34_5_, in1_34_6_, in1_34_7_, in1_34_8_, in1_34_9_,
     in1_34_10_, in1_34_11_, in1_34_24_, in1_35_0_, in1_35_1_, in1_35_2_,
     in1_35_3_, in1_35_4_, in1_35_5_, in1_35_6_, in1_35_7_, in1_35_8_, in1_35_9_,
     in1_35_10_, in1_35_11_, in1_37_0_, in1_37_1_, in1_37_2_, in1_37_3_,
     in1_37_4_, in1_37_5_, in1_37_6_, in1_37_7_, in1_37_8_, in1_37_9_,
     in1_37_10_, in1_37_11_, in1_37_12_, in1_37_24_, in1_38_0_, in1_38_1_,
     in1_38_2_, in1_38_3_, in1_38_4_, in1_38_5_, in1_38_6_, in1_38_7_, in1_38_8_,
     in1_38_9_, in1_38_10_, in1_38_11_, in1_38_12_, in1_40_0_, in1_40_1_,
     in1_40_2_, in1_40_3_, in1_40_4_, in1_40_5_, in1_40_6_, in1_40_7_, in1_40_8_,
     in1_40_9_, in1_40_10_, in1_40_11_, in1_40_12_, in1_40_13_, in1_40_24_,
     in1_41_0_, in1_41_1_, in1_41_2_, in1_41_3_, in1_41_4_, in1_41_5_, in1_41_6_,
     in1_41_7_, in1_41_8_, in1_41_9_, in1_41_10_, in1_41_11_, in1_41_12_,
     in1_41_13_, in1_43_0_, in1_43_1_, in1_43_2_, in1_43_3_, in1_43_4_,
     in1_43_5_, in1_43_6_, in1_43_7_, in1_43_8_, in1_43_9_, in1_43_10_,
     in1_43_11_, in1_43_12_, in1_43_13_, in1_43_14_, in1_43_24_, in1_44_0_,
     in1_44_1_, in1_44_2_, in1_44_3_, in1_44_4_, in1_44_5_, in1_44_6_, in1_44_7_,
     in1_44_8_, in1_44_9_, in1_44_10_, in1_44_11_, in1_44_12_, in1_44_13_,
     in1_44_14_, in1_46_0_, in1_46_1_, in1_46_2_, in1_46_3_, in1_46_4_,
     in1_46_5_, in1_46_6_, in1_46_7_, in1_46_8_, in1_46_9_, in1_46_10_,
     in1_46_11_, in1_46_12_, in1_46_13_, in1_46_14_, in1_46_15_, in1_46_24_,
     in1_47_0_, in1_47_1_, in1_47_2_, in1_47_3_, in1_47_4_, in1_47_5_, in1_47_6_,
     in1_47_7_, in1_47_8_, in1_47_9_, in1_47_10_, in1_47_11_, in1_47_12_,
     in1_47_13_, in1_47_14_, in1_47_15_, in1_49_0_, in1_49_1_, in1_49_2_,
     in1_49_3_, in1_49_4_, in1_49_5_, in1_49_6_, in1_49_7_, in1_49_8_, in1_49_9_,
     in1_49_10_, in1_49_11_, in1_49_12_, in1_49_13_, in1_49_14_, in1_49_15_,
     in1_49_16_, in1_49_24_, in1_50_0_, in1_50_1_, in1_50_2_, in1_50_3_,
     in1_50_4_, in1_50_5_, in1_50_6_, in1_50_7_, in1_50_8_, in1_50_9_,
     in1_50_10_, in1_50_11_, in1_50_12_, in1_50_13_, in1_50_14_, in1_50_15_,
     in1_50_16_, in1_52_0_, in1_52_1_, in1_52_2_, in1_52_3_, in1_52_4_,
     in1_52_5_, in1_52_6_, in1_52_7_, in1_52_8_, in1_52_9_, in1_52_10_,
     in1_52_11_, in1_52_12_, in1_52_13_, in1_52_14_, in1_52_15_, in1_52_16_,
     in1_52_17_, in1_52_24_, in1_53_0_, in1_53_1_, in1_53_2_, in1_53_3_,
     in1_53_4_, in1_53_5_, in1_53_6_, in1_53_7_, in1_53_8_, in1_53_9_,
     in1_53_10_, in1_53_11_, in1_53_12_, in1_53_13_, in1_53_14_, in1_53_15_,
     in1_53_16_, in1_53_17_, in1_55_0_, in1_55_1_, in1_55_2_, in1_55_3_,
     in1_55_4_, in1_55_5_, in1_55_6_, in1_55_7_, in1_55_8_, in1_55_9_,
     in1_55_10_, in1_55_11_, in1_55_12_, in1_55_13_, in1_55_14_, in1_55_15_,
     in1_55_16_, in1_55_17_, in1_55_18_, in1_55_24_, in1_56_0_, in1_56_1_,
     in1_56_2_, in1_56_3_, in1_56_4_, in1_56_5_, in1_56_6_, in1_56_7_, in1_56_8_,
     in1_56_9_, in1_56_10_, in1_56_11_, in1_56_12_, in1_56_13_, in1_56_14_,
     in1_56_15_, in1_56_16_, in1_56_17_, in1_56_18_, in1_58_0_, in1_58_1_,
     in1_58_2_, in1_58_3_, in1_58_4_, in1_58_5_, in1_58_6_, in1_58_7_, in1_58_8_,
     in1_58_9_, in1_58_10_, in1_58_11_, in1_58_12_, in1_58_13_, in1_58_14_,
     in1_58_15_, in1_58_16_, in1_58_17_, in1_58_18_, in1_58_19_, in1_58_24_,
     in1_59_0_, in1_59_1_, in1_59_2_, in1_59_3_, in1_59_4_, in1_59_5_, in1_59_6_,
     in1_59_7_, in1_59_8_, in1_59_9_, in1_59_10_, in1_59_11_, in1_59_12_,
     in1_59_13_, in1_59_14_, in1_59_15_, in1_59_16_, in1_59_17_, in1_59_18_,
     in1_59_19_, in1_61_0_, in1_61_1_, in1_61_2_, in1_61_3_, in1_61_4_,
     in1_61_5_, in1_61_6_, in1_61_7_, in1_61_8_, in1_61_9_, in1_61_10_,
     in1_61_11_, in1_61_12_, in1_61_13_, in1_61_14_, in1_61_15_, in1_61_16_,
     in1_61_17_, in1_61_18_, in1_61_19_, in1_61_20_, in1_61_24_, in1_62_0_,
     in1_62_1_, in1_62_2_, in1_62_3_, in1_62_4_, in1_62_5_, in1_62_6_, in1_62_7_,
     in1_62_8_, in1_62_9_, in1_62_10_, in1_62_11_, in1_62_12_, in1_62_13_,
     in1_62_14_, in1_62_15_, in1_62_16_, in1_62_17_, in1_62_18_, in1_62_19_,
     in1_62_20_, in1_64_0_, in1_64_1_, in1_64_2_, in1_64_3_, in1_64_4_,
     in1_64_5_, in1_64_6_, in1_64_7_, in1_64_8_, in1_64_9_, in1_64_10_,
     in1_64_11_, in1_64_12_, in1_64_13_, in1_64_14_, in1_64_15_, in1_64_16_,
     in1_64_17_, in1_64_18_, in1_64_19_, in1_64_20_, in1_64_21_, in1_64_24_,
     in1_65_0_, in1_65_1_, in1_65_2_, in1_65_3_, in1_65_4_, in1_65_5_, in1_65_6_,
     in1_65_7_, in1_65_8_, in1_65_9_, in1_65_10_, in1_65_11_, in1_65_12_,
     in1_65_13_, in1_65_14_, in1_65_15_, in1_65_16_, in1_65_17_, in1_65_18_,
     in1_65_19_, in1_65_20_, in1_65_21_, in1_67_0_, in1_67_1_, in1_67_2_,
     in1_67_3_, in1_67_4_, in1_67_5_, in1_67_6_, in1_67_7_, in1_67_8_, in1_67_9_,
     in1_67_10_, in1_67_11_, in1_67_12_, in1_67_13_, in1_67_14_, in1_67_15_,
     in1_67_16_, in1_67_17_, in1_67_18_, in1_67_19_, in1_67_20_, in1_67_21_,
     in1_67_22_, in1_67_24_, in1_68_0_, in1_68_1_, in1_68_2_, in1_68_3_,
     in1_68_4_, in1_68_5_, in1_68_6_, in1_68_7_, in1_68_8_, in1_68_9_,
     in1_68_10_, in1_68_11_, in1_68_12_, in1_68_13_, in1_68_14_, in1_68_15_,
     in1_68_16_, in1_68_17_, in1_68_18_, in1_68_19_, in1_68_20_, in1_68_21_,
     in1_68_22_, in1_70_0_, in1_70_1_, in1_70_2_, in1_70_3_, in1_70_4_,
     in1_70_5_, in1_70_6_, in1_70_7_, in1_70_8_, in1_70_9_, in1_70_10_,
     in1_70_11_, in1_70_12_, in1_70_13_, in1_70_14_, in1_70_15_, in1_70_16_,
     in1_70_17_, in1_70_18_, in1_70_19_, in1_70_20_, in1_70_21_, in1_70_22_,
     in1_70_23_, in1_70_24_, in1_71_0_, in1_71_1_, in1_71_2_, in1_71_3_,
     in1_71_4_, in1_71_5_, in1_71_6_, in1_71_7_, in1_71_8_, in1_71_9_,
     in1_71_10_, in1_71_11_, in1_71_12_, in1_71_13_, in1_71_14_, in1_71_15_,
     in1_71_16_, in1_71_17_, in1_71_18_, in1_71_19_, in1_71_20_, in1_71_21_,
     in1_71_22_, in1_71_23_, in1_73_0_, in1_73_1_, in1_73_2_, in1_73_3_,
     in1_73_4_, in1_73_5_, in1_73_6_, in1_73_7_, in1_73_8_, in1_73_9_,
     in1_73_10_, in1_73_11_, in1_73_12_, in1_73_13_, in1_73_14_, in1_73_15_,
     in1_73_16_, in1_73_17_, in1_73_18_, in1_73_19_, in1_73_20_, in1_73_21_,
     in1_73_22_, in1_73_23_, in1_73_24_, in1_74_0_, in1_74_1_, in1_74_2_,
     in1_74_3_, in1_74_4_, in1_74_5_, in1_74_6_, in1_74_7_, in1_74_8_, in1_74_9_,
     in1_74_10_, in1_74_11_, in1_74_12_, in1_74_13_, in1_74_14_, in1_74_15_,
     in1_74_16_, in1_74_17_, in1_74_18_, in1_74_19_, in1_74_20_, in1_74_21_,
     in1_74_22_, in1_74_23_, in1_76_0_, in1_76_1_, in1_76_2_, in1_76_3_,
     in1_76_4_, in1_76_5_, in1_76_6_, in1_76_7_, in1_76_8_, in1_76_9_,
     in1_76_10_, in1_76_11_, in1_76_12_, in1_76_13_, in1_76_14_, in1_76_15_,
     in1_76_16_, in1_76_17_, in1_76_18_, in1_76_19_, in1_76_20_, in1_76_21_,
     in1_76_22_, in1_76_23_, in1_76_24_, in1_77_0_, in1_77_1_, in1_77_2_,
     in1_77_3_, in1_77_4_, in1_77_5_, in1_77_6_, in1_77_7_, in1_77_8_, in1_77_9_,
     in1_77_10_, in1_77_11_, in1_77_12_, in1_77_13_, in1_77_14_, in1_77_15_,
     in1_77_16_, in1_77_17_, in1_77_18_, in1_77_19_, in1_77_20_, in1_77_21_,
     in1_77_22_, in1_77_23_, in1_79_0_, in1_79_1_, in1_79_2_, in1_79_3_,
     in1_79_4_, in1_79_5_, in1_79_6_, in1_79_7_, in1_79_8_, in1_79_9_,
     in1_79_10_, in1_79_11_, in1_79_12_, in1_79_13_, in1_79_14_, in1_79_15_,
     in1_79_16_, in1_79_17_, in1_79_18_, in1_79_19_, in1_79_20_, in1_79_21_,
     in1_79_22_, in1_79_23_, in1_79_24_, in1_80_0_, in1_80_1_, in1_80_2_,
     in1_80_3_, in1_80_4_, in1_80_5_, in1_80_6_, in1_80_7_, in1_80_8_, in1_80_9_,
     in1_80_10_, in1_80_11_, in1_80_12_, in1_80_13_, in1_80_14_, in1_80_15_,
     in1_80_16_, in1_80_17_, in1_80_18_, in1_80_19_, in1_80_20_, in1_80_21_,
     in1_80_22_, in1_80_23_, in1_82_0_, in1_82_1_, in1_82_2_, in1_82_3_,
     in1_82_4_, in1_82_5_, in1_82_6_, in1_82_7_, in1_82_8_, in1_82_9_,
     in1_82_10_, in1_82_11_, in1_82_12_, in1_82_13_, in1_82_14_, in1_82_15_,
     in1_82_16_, in1_82_17_, in1_82_18_, in1_82_19_, in1_82_20_, in1_82_21_,
     in1_82_22_, in1_82_23_, in1_82_24_, in1_83_0_, in1_83_1_, in1_83_2_,
     in1_83_3_, in1_83_4_, in1_83_5_, in1_83_6_, in1_83_7_, in1_83_8_, in1_83_9_,
     in1_83_10_, in1_83_11_, in1_83_12_, in1_83_13_, in1_83_14_, in1_83_15_,
     in1_83_16_, in1_83_17_, in1_83_18_, in1_83_19_, in1_83_20_, in1_83_21_,
     in1_83_22_, in1_83_23_, in1_85_0_, in1_85_1_, in1_85_2_, in1_85_3_,
     in1_85_4_, in1_85_5_, in1_85_6_, in1_85_7_, in1_85_8_, in1_85_9_,
     in1_85_10_, in1_85_11_, in1_85_12_, in1_85_13_, in1_85_14_, in1_85_15_,
     in1_85_16_, in1_85_17_, in1_85_18_, in1_85_19_, in1_85_20_, in1_85_21_,
     in1_85_22_, in1_85_23_, in1_85_24_, in1_86_0_, in1_86_1_, in1_86_2_,
     in1_86_3_, in1_86_4_, in1_86_5_, in1_86_6_, in1_86_7_, in1_86_8_, in1_86_9_,
     in1_86_10_, in1_86_11_, in1_86_12_, in1_86_13_, in1_86_14_, in1_86_15_,
     in1_86_16_, in1_86_17_, in1_86_18_, in1_86_19_, in1_86_20_, in1_86_21_,
     in1_86_22_, in1_86_23_, in1_88_0_, in1_88_1_, in1_88_2_, in1_88_3_,
     in1_88_4_, in1_88_5_, in1_88_6_, in1_88_7_, in1_88_8_, in1_88_9_,
     in1_88_10_, in1_88_11_, in1_88_12_, in1_88_13_, in1_88_14_, in1_88_15_,
     in1_88_16_, in1_88_17_, in1_88_18_, in1_88_19_, in1_88_20_, in1_88_21_,
     in1_88_22_, in1_88_23_, in1_88_24_, in1_89_0_, in1_89_1_, in1_89_2_,
     in1_89_3_, in1_89_4_, in1_89_5_, in1_89_6_, in1_89_7_, in1_89_8_, in1_89_9_,
     in1_89_10_, in1_89_11_, in1_89_12_, in1_89_13_, in1_89_14_, in1_89_15_,
     in1_89_16_, in1_89_17_, in1_89_18_, in1_89_19_, in1_89_20_, in1_89_21_,
     in1_89_22_, in1_89_23_, in1_91_0_, in1_91_1_, in1_91_2_, in1_91_3_,
     in1_91_4_, in1_91_5_, in1_91_6_, in1_91_7_, in1_91_8_, in1_91_9_,
     in1_91_10_, in1_91_11_, in1_91_12_, in1_91_13_, in1_91_14_, in1_91_15_,
     in1_91_16_, in1_91_17_, in1_91_18_, in1_91_19_, in1_91_20_, in1_91_21_,
     in1_91_22_, in1_91_23_, in1_91_24_, in1_92_0_, in1_92_1_, in1_92_2_,
     in1_92_3_, in1_92_4_, in1_92_5_, in1_92_6_, in1_92_7_, in1_92_8_, in1_92_9_,
     in1_92_10_, in1_92_11_, in1_92_12_, in1_92_13_, in1_92_14_, in1_92_15_,
     in1_92_16_, in1_92_17_, in1_92_18_, in1_92_19_, in1_92_20_, in1_92_21_,
     in1_92_22_, in1_92_23_, in1_94_0_, in1_94_1_, in1_94_2_, in1_94_3_,
     in1_94_4_, in1_94_5_, in1_94_6_, in1_94_7_, in1_94_8_, in1_94_9_,
     in1_94_10_, in1_94_11_, in1_94_12_, in1_94_13_, in1_94_14_, in1_94_15_,
     in1_94_16_, in1_94_17_, in1_94_18_, in1_94_19_, in1_94_20_, in1_94_21_,
     in1_94_22_, in1_94_23_, in1_94_24_, in1_95_0_, in1_95_1_, in1_95_2_,
     in1_95_3_, in1_95_4_, in1_95_5_, in1_95_6_, in1_95_7_, in1_95_8_, in1_95_9_,
     in1_95_10_, in1_95_11_, in1_95_12_, in1_95_13_, in1_95_14_, in1_95_15_,
     in1_95_16_, in1_95_17_, in1_95_18_, in1_95_19_, in1_95_20_, in1_95_21_,
     in1_95_22_, in1_95_23_, in1_97_0_, in1_97_1_, in1_97_2_, in1_97_3_,
     in1_97_4_, in1_97_5_, in1_97_6_, in1_97_7_, in1_97_8_, in1_97_9_,
     in1_97_10_, in1_97_11_, in1_97_12_, in1_97_13_, in1_97_14_, in1_97_15_,
     in1_97_16_, in1_97_17_, in1_97_18_, in1_97_19_, in1_97_20_, in1_97_21_,
     in1_97_22_, in1_97_23_, in1_97_24_, in1_98_0_, in1_98_1_, in1_98_2_,
     in1_98_3_, in1_98_4_, in1_98_5_, in1_98_6_, in1_98_7_, in1_98_8_, in1_98_9_,
     in1_98_10_, in1_98_11_, in1_98_12_, in1_98_13_, in1_98_14_, in1_98_15_,
     in1_98_16_, in1_98_17_, in1_98_18_, in1_98_19_, in1_98_20_, in1_98_21_,
     in1_98_22_, in1_98_23_, in1_100_0_, in1_100_1_, in1_100_2_, in1_100_3_,
     in1_100_4_, in1_100_5_, in1_100_6_, in1_100_7_, in1_100_8_, in1_100_9_,
     in1_100_10_, in1_100_11_, in1_100_12_, in1_100_13_, in1_100_14_,
     in1_100_15_, in1_100_16_, in1_100_17_, in1_100_18_, in1_100_19_,
     in1_100_20_, in1_100_21_, in1_100_22_, in1_100_23_, in1_100_24_, in1_101_0_,
     in1_101_1_, in1_101_2_, in1_101_3_, in1_101_4_, in1_101_5_, in1_101_6_,
     in1_101_7_, in1_101_8_, in1_101_9_, in1_101_10_, in1_101_11_, in1_101_12_,
     in1_101_13_, in1_101_14_, in1_101_15_, in1_101_16_, in1_101_17_,
     in1_101_18_, in1_101_19_, in1_101_20_, in1_101_21_, in1_101_22_,
     in1_101_23_, in1_103_0_, in1_103_1_, in1_103_2_, in1_103_3_, in1_103_4_,
     in1_103_5_, in1_103_6_, in1_103_7_, in1_103_8_, in1_103_9_, in1_103_10_,
     in1_103_11_, in1_103_12_, in1_103_13_, in1_103_14_, in1_103_15_,
     in1_103_16_, in1_103_17_, in1_103_18_, in1_103_19_, in1_103_20_,
     in1_103_21_, in1_103_22_, in1_103_23_, in1_103_24_, in1_104_0_, in1_104_1_,
     in1_104_2_, in1_104_3_, in1_104_4_, in1_104_5_, in1_104_6_, in1_104_7_,
     in1_104_8_, in1_104_9_, in1_104_10_, in1_104_11_, in1_104_12_, in1_104_13_,
     in1_104_14_, in1_104_15_, in1_104_16_, in1_104_17_, in1_104_18_,
     in1_104_19_, in1_104_20_, in1_104_21_, in1_104_22_, in1_104_23_, in1_106_0_,
     in1_106_1_, in1_106_2_, in1_106_3_, in1_106_4_, in1_106_5_, in1_106_6_,
     in1_106_7_, in1_106_8_, in1_106_9_, in1_106_10_, in1_106_11_, in1_106_12_,
     in1_106_13_, in1_106_14_, in1_106_15_, in1_106_16_, in1_106_17_,
     in1_106_18_, in1_106_19_, in1_106_20_, in1_106_21_, in1_106_22_,
     in1_106_23_, in1_106_24_, in1_107_0_, in1_107_1_, in1_107_2_, in1_107_3_,
     in1_107_4_, in1_107_5_, in1_107_6_, in1_107_7_, in1_107_8_, in1_107_9_,
     in1_107_10_, in1_107_11_, in1_107_12_, in1_107_13_, in1_107_14_,
     in1_107_15_, in1_107_16_, in1_107_17_, in1_107_18_, in1_107_19_,
     in1_107_20_, in1_107_21_, in1_107_22_, in1_107_23_, in1_109_0_, in1_109_1_,
     in1_109_2_, in1_109_3_, in1_109_4_, in1_109_5_, in1_109_6_, in1_109_7_,
     in1_109_8_, in1_109_9_, in1_109_10_, in1_109_11_, in1_109_12_, in1_109_13_,
     in1_109_14_, in1_109_15_, in1_109_16_, in1_109_17_, in1_109_18_,
     in1_109_19_, in1_109_20_, in1_109_21_, in1_109_22_, in1_109_23_,
     in1_109_24_, in1_110_0_, in1_110_1_, in1_110_2_, in1_110_3_, in1_110_4_,
     in1_110_5_, in1_110_6_, in1_110_7_, in1_110_8_, in1_110_9_, in1_110_10_,
     in1_110_11_, in1_110_12_, in1_110_13_, in1_110_14_, in1_110_15_,
     in1_110_16_, in1_110_17_, in1_110_18_, in1_110_19_, in1_110_20_,
     in1_110_21_, in1_110_22_, in1_110_23_, in1_112_0_, in1_112_1_, in1_112_2_,
     in1_112_3_, in1_112_4_, in1_112_5_, in1_112_6_, in1_112_7_, in1_112_8_,
     in1_112_9_, in1_112_10_, in1_112_11_, in1_112_12_, in1_112_13_, in1_112_14_,
     in1_112_15_, in1_112_16_, in1_112_17_, in1_112_18_, in1_112_19_,
     in1_112_20_, in1_112_21_, in1_112_22_, in1_112_23_, in1_112_24_, in1_113_0_,
     in1_113_1_, in1_113_2_, in1_113_3_, in1_113_4_, in1_113_5_, in1_113_6_,
     in1_113_7_, in1_113_8_, in1_113_9_, in1_113_10_, in1_113_11_, in1_113_12_,
     in1_113_13_, in1_113_14_, in1_113_15_, in1_113_16_, in1_113_17_,
     in1_113_18_, in1_113_19_, in1_113_20_, in1_113_21_, in1_113_22_,
     in1_113_23_, in1_115_0_, in1_115_1_, in1_115_2_, in1_115_3_, in1_115_4_,
     in1_115_5_, in1_115_6_, in1_115_7_, in1_115_8_, in1_115_9_, in1_115_10_,
     in1_115_11_, in1_115_12_, in1_115_13_, in1_115_14_, in1_115_15_,
     in1_115_16_, in1_115_17_, in1_115_18_, in1_115_19_, in1_115_20_,
     in1_115_21_, in1_115_22_, in1_115_23_, in1_115_24_, in1_116_0_, in1_116_1_,
     in1_116_2_, in1_116_3_, in1_116_4_, in1_116_5_, in1_116_6_, in1_116_7_,
     in1_116_8_, in1_116_9_, in1_116_10_, in1_116_11_, in1_116_12_, in1_116_13_,
     in1_116_14_, in1_116_15_, in1_116_16_, in1_116_17_, in1_116_18_,
     in1_116_19_, in1_116_20_, in1_116_21_, in1_116_22_, in1_116_23_, in1_118_0_,
     in1_118_1_, in1_118_2_, in1_118_3_, in1_118_4_, in1_118_5_, in1_118_6_,
     in1_118_7_, in1_118_8_, in1_118_9_, in1_118_10_, in1_118_11_, in1_118_12_,
     in1_118_13_, in1_118_14_, in1_118_15_, in1_118_16_, in1_118_17_,
     in1_118_18_, in1_118_19_, in1_118_20_, in1_118_21_, in1_118_22_,
     in1_118_23_, in1_118_24_, in1_119_0_, in1_119_1_, in1_119_2_, in1_119_3_,
     in1_119_4_, in1_119_5_, in1_119_6_, in1_119_7_, in1_119_8_, in1_119_9_,
     in1_119_10_, in1_119_11_, in1_119_12_, in1_119_13_, in1_119_14_,
     in1_119_15_, in1_119_16_, in1_119_17_, in1_119_18_, in1_119_19_,
     in1_119_20_, in1_119_21_, in1_119_22_, in1_119_23_, in1_121_0_, in1_121_1_,
     in1_121_2_, in1_121_3_, in1_121_4_, in1_121_5_, in1_121_6_, in1_121_7_,
     in1_121_8_, in1_121_9_, in1_121_10_, in1_121_11_, in1_121_12_, in1_121_13_,
     in1_121_14_, in1_121_15_, in1_121_16_, in1_121_17_, in1_121_18_,
     in1_121_19_, in1_121_20_, in1_121_21_, in1_121_22_, in1_121_23_,
     in1_121_24_, in1_122_0_, in1_122_1_, in1_122_2_, in1_122_3_, in1_122_4_,
     in1_122_5_, in1_122_6_, in1_122_7_, in1_122_8_, in1_122_9_, in1_122_10_,
     in1_122_11_, in1_122_12_, in1_122_13_, in1_122_14_, in1_122_15_,
     in1_122_16_, in1_122_17_, in1_122_18_, in1_122_19_, in1_122_20_,
     in1_122_21_, in1_122_22_, in1_122_23_, in1_124_0_, in1_124_1_, in1_124_2_,
     in1_124_3_, in1_124_4_, in1_124_5_, in1_124_6_, in1_124_7_, in1_124_8_,
     in1_124_9_, in1_124_10_, in1_124_11_, in1_124_12_, in1_124_13_, in1_124_14_,
     in1_124_15_, in1_124_16_, in1_124_17_, in1_124_18_, in1_124_19_,
     in1_124_20_, in1_124_21_, in1_124_22_, in1_124_23_, in1_124_24_, in1_125_0_,
     in1_125_1_, in1_125_2_, in1_125_3_, in1_125_4_, in1_125_5_, in1_125_6_,
     in1_125_7_, in1_125_8_, in1_125_9_, in1_125_10_, in1_125_11_, in1_125_12_,
     in1_125_13_, in1_125_14_, in1_125_15_, in1_125_16_, in1_125_17_,
     in1_125_18_, in1_125_19_, in1_125_20_, in1_125_21_, in1_125_22_,
     in1_125_23_, in1_127_0_, in1_127_1_, in1_127_2_, in1_127_3_, in1_127_4_,
     in1_127_5_, in1_127_6_, in1_127_7_, in1_127_8_, in1_127_9_, in1_127_10_,
     in1_127_11_, in1_127_12_, in1_127_13_, in1_127_14_, in1_127_15_,
     in1_127_16_, in1_127_17_, in1_127_18_, in1_127_19_, in1_127_20_,
     in1_127_21_, in1_127_22_, in1_127_23_, in1_127_24_, in1_128_0_, in1_128_1_,
     in1_128_2_, in1_128_3_, in1_128_4_, in1_128_5_, in1_128_6_, in1_128_7_,
     in1_128_8_, in1_128_9_, in1_128_10_, in1_128_11_, in1_128_12_, in1_128_13_,
     in1_128_14_, in1_128_15_, in1_128_16_, in1_128_17_, in1_128_18_,
     in1_128_19_, in1_128_20_, in1_128_21_, in1_128_22_, in1_128_23_, in1_130_0_,
     in1_130_1_, in1_130_2_, in1_130_3_, in1_130_4_, in1_130_5_, in1_130_6_,
     in1_130_7_, in1_130_8_, in1_130_9_, in1_130_10_, in1_130_11_, in1_130_12_,
     in1_130_13_, in1_130_14_, in1_130_15_, in1_130_16_, in1_130_17_,
     in1_130_18_, in1_130_19_, in1_130_20_, in1_130_21_, in1_130_22_,
     in1_130_23_, in1_130_24_, in1_131_0_, in1_131_1_, in1_131_2_, in1_131_3_,
     in1_131_4_, in1_131_5_, in1_131_6_, in1_131_7_, in1_131_8_, in1_131_9_,
     in1_131_10_, in1_131_11_, in1_131_12_, in1_131_13_, in1_131_14_,
     in1_131_15_, in1_131_16_, in1_131_17_, in1_131_18_, in1_131_19_,
     in1_131_20_, in1_131_21_, in1_131_22_, in1_131_23_, in1_133_0_, in1_133_1_,
     in1_133_2_, in1_133_3_, in1_133_4_, in1_133_5_, in1_133_6_, in1_133_7_,
     in1_133_8_, in1_133_9_, in1_133_10_, in1_133_11_, in1_133_12_, in1_133_13_,
     in1_133_14_, in1_133_15_, in1_133_16_, in1_133_17_, in1_133_18_,
     in1_133_19_, in1_133_20_, in1_133_21_, in1_133_22_, in1_133_23_,
     in1_133_24_, in1_134_0_, in1_134_1_, in1_134_2_, in1_134_3_, in1_134_4_,
     in1_134_5_, in1_134_6_, in1_134_7_, in1_134_8_, in1_134_9_, in1_134_10_,
     in1_134_11_, in1_134_12_, in1_134_13_, in1_134_14_, in1_134_15_,
     in1_134_16_, in1_134_17_, in1_134_18_, in1_134_19_, in1_134_20_,
     in1_134_21_, in1_134_22_, in1_134_23_, in1_136_0_, in1_136_1_, in1_136_2_,
     in1_136_3_, in1_136_4_, in1_136_5_, in1_136_6_, in1_136_7_, in1_136_8_,
     in1_136_9_, in1_136_10_, in1_136_11_, in1_136_12_, in1_136_13_, in1_136_14_,
     in1_136_15_, in1_136_16_, in1_136_17_, in1_136_18_, in1_136_19_,
     in1_136_20_, in1_136_21_, in1_136_22_, in1_136_23_, in1_136_24_, in1_137_0_,
     in1_137_1_, in1_137_2_, in1_137_3_, in1_137_4_, in1_137_5_, in1_137_6_,
     in1_137_7_, in1_137_8_, in1_137_9_, in1_137_10_, in1_137_11_, in1_137_12_,
     in1_137_13_, in1_137_14_, in1_137_15_, in1_137_16_, in1_137_17_,
     in1_137_18_, in1_137_19_, in1_137_20_, in1_137_21_, in1_137_22_,
     in1_137_23_, in1_139_0_, in1_139_1_, in1_139_2_, in1_139_3_, in1_139_4_,
     in1_139_5_, in1_139_6_, in1_139_7_, in1_139_8_, in1_139_9_, in1_139_10_,
     in1_139_11_, in1_139_12_, in1_139_13_, in1_139_14_, in1_139_15_,
     in1_139_16_, in1_139_17_, in1_139_18_, in1_139_19_, in1_139_20_,
     in1_139_21_, in1_139_22_, in1_139_23_, in1_139_24_, in1_140_0_, in1_140_1_,
     in1_140_2_, in1_140_3_, in1_140_4_, in1_140_5_, in1_140_6_, in1_140_7_,
     in1_140_8_, in1_140_9_, in1_140_10_, in1_140_11_, in1_140_12_, in1_140_13_,
     in1_140_14_, in1_140_15_, in1_140_16_, in1_140_17_, in1_140_18_,
     in1_140_19_, in1_140_20_, in1_140_21_, in1_140_22_, in1_140_23_, in1_142_0_,
     in1_142_1_, in1_142_2_, in1_142_3_, in1_142_4_, in1_142_5_, in1_142_6_,
     in1_142_7_, in1_142_8_, in1_142_9_, in1_142_10_, in1_142_11_, in1_142_12_,
     in1_142_13_, in1_142_14_, in1_142_15_, in1_142_16_, in1_142_17_,
     in1_142_18_, in1_142_19_, in1_142_20_, in1_142_21_, in1_142_22_,
     in1_142_23_, in1_142_24_, in1_143_0_, in1_143_1_, in1_143_2_, in1_143_3_,
     in1_143_4_, in1_143_5_, in1_143_6_, in1_143_7_, in1_143_8_, in1_143_9_,
     in1_143_10_, in1_143_11_, in1_143_12_, in1_143_13_, in1_143_14_,
     in1_143_15_, in1_143_16_, in1_143_17_, in1_143_18_, in1_143_19_,
     in1_143_20_, in1_143_21_, in1_143_22_, in1_143_23_, in1_145_24_;
assign n_1285 = asc001_0_36_;
assign n_1286 = asc001_0_35_;
assign n_1287 = asc001_0_34_;
assign n_1288 = asc001_0_33_;
assign n_1289 = asc001_0_32_;
assign n_1290 = asc001_0_31_;
assign n_1291 = asc001_0_30_;
assign n_1292 = asc001_0_29_;
assign n_1293 = asc001_0_28_;
assign n_1294 = asc001_0_27_;
assign n_1295 = asc001_0_26_;
assign n_1296 = asc001_0_25_;
assign n_1297 = asc001_0_24_;
assign n_1298 = asc001_0_23_;
assign n_1299 = asc001_0_22_;
assign n_1300 = asc001_0_21_;
assign n_1301 = asc001_0_20_;
assign n_1302 = asc001_0_19_;
assign n_1303 = asc001_0_18_;
assign n_1304 = asc001_0_17_;
assign n_1305 = asc001_0_16_;
assign n_1306 = asc001_0_15_;
assign n_1307 = asc001_0_14_;
assign n_1308 = asc001_0_13_;
assign n_1309 = asc001_0_12_;
assign n_1310 = asc001_0_11_;
assign n_1311 = asc001_0_10_;
assign n_1312 = asc001_0_9_;
assign n_1313 = asc001_0_8_;
assign n_1314 = asc001_0_7_;
assign n_1315 = asc001_0_6_;
assign n_1316 = asc001_0_5_;
assign n_1317 = asc001_0_4_;
assign n_1318 = asc001_0_3_;
assign n_1319 = asc001_0_2_;
assign n_1320 = asc001_0_1_;
assign n_1321 = asc001_0_0_;
assign {out1[34]} = n_1287;
assign {out1[32]} = n_1289;
assign {out1[29]} = n_1292;
assign {out1[28]} = n_1293;
assign {out1[23]} = n_1298;
assign {out1[21]} = n_1300;
assign {out1[20]} = n_1301;
assign {out1[19]} = n_1302;
assign {out1[18]} = n_1303;
assign {out1[17]} = n_1304;
assign {out1[16]} = n_1305;
assign {out1[15]} = n_1306;
assign {out1[14]} = n_1307;
assign {out1[13]} = n_1308;
assign {out1[12]} = n_1309;
assign {out1[11]} = n_1310;
assign {out1[10]} = n_1311;
assign {out1[9]} = n_1312;
assign {out1[8]} = n_1313;
assign {out1[7]} = n_1314;
assign {out1[6]} = n_1315;
assign {out1[5]} = n_1316;
assign {out1[4]} = n_1317;
assign {out1[3]} = n_1318;
assign {out1[2]} = n_1319;
assign {out1[1]} = n_1320;
assign {out1[0]} = n_1321;
reg cadence_register_n_1397;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1397 <= in1[0];
    end
 end
 assign n_1397 = cadence_register_n_1397;
reg cadence_register_n_1398;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1398 <= n_1397;
    end
 end
 assign n_1398 = cadence_register_n_1398;
reg cadence_register_n_1399;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1399 <= in1[1];
    end
 end
 assign n_1399 = cadence_register_n_1399;
reg cadence_register_n_1400;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1400 <= n_1399;
    end
 end
 assign n_1400 = cadence_register_n_1400;
reg cadence_register_n_1401;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1401 <= in1[8];
    end
 end
 assign n_1401 = cadence_register_n_1401;
reg cadence_register_n_1402;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1402 <= n_1401;
    end
 end
 assign n_1402 = cadence_register_n_1402;
reg cadence_register_n_1403;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1403 <= in2[23];
    end
 end
 assign n_1403 = cadence_register_n_1403;
reg cadence_register_n_1404;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1404 <= n_1403;
    end
 end
 assign n_1404 = cadence_register_n_1404;
reg cadence_register_n_1405;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1405 <= sub_949_2_n_76;
    end
 end
 assign n_1405 = cadence_register_n_1405;
reg cadence_register_n_1406;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1406 <= in1_85_24_;
    end
 end
 assign n_1406 = cadence_register_n_1406;
reg cadence_register_n_1407;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1407 <= in1_100_24_;
    end
 end
 assign n_1407 = cadence_register_n_1407;
reg cadence_register_n_1408;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1408 <= in1_88_24_;
    end
 end
 assign n_1408 = cadence_register_n_1408;
reg cadence_register_n_1409;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1409 <= in1_107_7_;
    end
 end
 assign n_1409 = cadence_register_n_1409;
reg cadence_register_n_1410;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1410 <= in1_107_5_;
    end
 end
 assign n_1410 = cadence_register_n_1410;
reg cadence_register_n_1411;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1411 <= in1_107_11_;
    end
 end
 assign n_1411 = cadence_register_n_1411;
reg cadence_register_n_1412;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1412 <= in1_109_13_;
    end
 end
 assign n_1412 = cadence_register_n_1412;
reg cadence_register_n_1413;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1413 <= in1_97_24_;
    end
 end
 assign n_1413 = cadence_register_n_1413;
reg cadence_register_n_1414;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1414 <= in1_94_24_;
    end
 end
 assign n_1414 = cadence_register_n_1414;
reg cadence_register_n_1415;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1415 <= in1_91_24_;
    end
 end
 assign n_1415 = cadence_register_n_1415;
reg cadence_register_n_1416;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1416 <= in1_109_12_;
    end
 end
 assign n_1416 = cadence_register_n_1416;
reg cadence_register_n_1417;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1417 <= sub_949_2_n_136;
    end
 end
 assign n_1417 = cadence_register_n_1417;
reg cadence_register_n_1418;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1418 <= sub_949_2_n_162;
    end
 end
 assign n_1418 = cadence_register_n_1418;
reg cadence_register_n_1419;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1419 <= sub_949_2_n_164;
    end
 end
 assign n_1419 = cadence_register_n_1419;
reg cadence_register_n_1420;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1420 <= in1_107_10_;
    end
 end
 assign n_1420 = cadence_register_n_1420;
reg cadence_register_n_1421;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1421 <= in1_107_15_;
    end
 end
 assign n_1421 = cadence_register_n_1421;
reg cadence_register_n_1422;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1422 <= in1_107_14_;
    end
 end
 assign n_1422 = cadence_register_n_1422;
reg cadence_register_n_1423;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1423 <= sub_949_2_n_12;
    end
 end
 assign n_1423 = cadence_register_n_1423;
reg cadence_register_n_1424;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1424 <= sub_949_2_n_147;
    end
 end
 assign n_1424 = cadence_register_n_1424;
reg cadence_register_n_1425;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1425 <= in1_107_4_;
    end
 end
 assign n_1425 = cadence_register_n_1425;
reg cadence_register_n_1426;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1426 <= in1_109_8_;
    end
 end
 assign n_1426 = cadence_register_n_1426;
reg cadence_register_n_1427;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1427 <= in1_109_6_;
    end
 end
 assign n_1427 = cadence_register_n_1427;
reg cadence_register_n_1428;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1428 <= in1_109_5_;
    end
 end
 assign n_1428 = cadence_register_n_1428;
reg cadence_register_n_1429;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1429 <= in1_109_10_;
    end
 end
 assign n_1429 = cadence_register_n_1429;
reg cadence_register_n_1430;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1430 <= in1_109_11_;
    end
 end
 assign n_1430 = cadence_register_n_1430;
reg cadence_register_n_1431;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1431 <= in1_107_3_;
    end
 end
 assign n_1431 = cadence_register_n_1431;
reg cadence_register_n_1432;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1432 <= in1_109_4_;
    end
 end
 assign n_1432 = cadence_register_n_1432;
reg cadence_register_n_1433;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1433 <= in1_107_2_;
    end
 end
 assign n_1433 = cadence_register_n_1433;
reg cadence_register_n_1434;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1434 <= in1_109_3_;
    end
 end
 assign n_1434 = cadence_register_n_1434;
reg cadence_register_n_1435;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1435 <= in1_107_12_;
    end
 end
 assign n_1435 = cadence_register_n_1435;
reg cadence_register_n_1436;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1436 <= in1_107_13_;
    end
 end
 assign n_1436 = cadence_register_n_1436;
reg cadence_register_n_1437;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1437 <= sub_949_2_n_7;
    end
 end
 assign n_1437 = cadence_register_n_1437;
reg cadence_register_n_1438;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1438 <= in1_103_24_;
    end
 end
 assign n_1438 = cadence_register_n_1438;
reg cadence_register_n_1439;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1439 <= in1_107_22_;
    end
 end
 assign n_1439 = cadence_register_n_1439;
reg cadence_register_n_1440;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1440 <= in1_106_24_;
    end
 end
 assign n_1440 = cadence_register_n_1440;
reg cadence_register_n_1441;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1441 <= in1_107_18_;
    end
 end
 assign n_1441 = cadence_register_n_1441;
reg cadence_register_n_1442;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1442 <= in1_107_21_;
    end
 end
 assign n_1442 = cadence_register_n_1442;
reg cadence_register_n_1443;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1443 <= in1_107_9_;
    end
 end
 assign n_1443 = cadence_register_n_1443;
reg cadence_register_n_1444;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1444 <= in1_107_20_;
    end
 end
 assign n_1444 = cadence_register_n_1444;
reg cadence_register_n_1445;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1445 <= in1_107_17_;
    end
 end
 assign n_1445 = cadence_register_n_1445;
reg cadence_register_n_1446;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1446 <= sub_949_2_n_50;
    end
 end
 assign n_1446 = cadence_register_n_1446;
reg cadence_register_n_1447;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1447 <= sub_949_2_n_51;
    end
 end
 assign n_1447 = cadence_register_n_1447;
reg cadence_register_n_1448;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1448 <= in1_107_1_;
    end
 end
 assign n_1448 = cadence_register_n_1448;
reg cadence_register_n_1449;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1449 <= in1_109_2_;
    end
 end
 assign n_1449 = cadence_register_n_1449;
reg cadence_register_n_1450;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1450 <= in1_107_19_;
    end
 end
 assign n_1450 = cadence_register_n_1450;
reg cadence_register_n_1451;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1451 <= in1_107_8_;
    end
 end
 assign n_1451 = cadence_register_n_1451;
reg cadence_register_n_1452;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1452 <= in1_109_9_;
    end
 end
 assign n_1452 = cadence_register_n_1452;
reg cadence_register_n_1453;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1453 <= sub_949_2_n_49;
    end
 end
 assign n_1453 = cadence_register_n_1453;
reg cadence_register_n_1454;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1454 <= in1_109_7_;
    end
 end
 assign n_1454 = cadence_register_n_1454;
reg cadence_register_n_1455;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1455 <= in1_107_6_;
    end
 end
 assign n_1455 = cadence_register_n_1455;
reg cadence_register_n_1456;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1456 <= in1_107_16_;
    end
 end
 assign n_1456 = cadence_register_n_1456;
reg cadence_register_n_1457;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1457 <= sub_949_2_n_63;
    end
 end
 assign n_1457 = cadence_register_n_1457;
reg cadence_register_n_1458;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1458 <= sub_949_2_n_55;
    end
 end
 assign n_1458 = cadence_register_n_1458;
reg cadence_register_n_1459;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1459 <= in1_107_23_;
    end
 end
 assign n_1459 = cadence_register_n_1459;
reg cadence_register_out1_26;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_26 <= n_1295;
    end
 end
 assign out1[26] = cadence_register_out1_26;
reg cadence_register_n_1461;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1461 <= in1_76_24_;
    end
 end
 assign n_1461 = cadence_register_n_1461;
reg cadence_register_n_1462;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1462 <= in1_82_24_;
    end
 end
 assign n_1462 = cadence_register_n_1462;
reg cadence_register_out1_22;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_22 <= n_1299;
    end
 end
 assign out1[22] = cadence_register_out1_22;
reg cadence_register_out1_24;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_24 <= n_1297;
    end
 end
 assign out1[24] = cadence_register_out1_24;
reg cadence_register_out1_25;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_25 <= n_1296;
    end
 end
 assign out1[25] = cadence_register_out1_25;
reg cadence_register_n_1466;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1466 <= sub_949_2_n_82;
    end
 end
 assign n_1466 = cadence_register_n_1466;
reg cadence_register_n_1467;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1467 <= in1_107_0_;
    end
 end
 assign n_1467 = cadence_register_n_1467;
reg cadence_register_n_1468;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1468 <= n_1286;
    end
 end
 assign n_1468 = cadence_register_n_1468;
reg cadence_register_out1_35;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_35 <= n_1468;
    end
 end
 assign out1[35] = cadence_register_out1_35;
reg cadence_register_n_1470;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1470 <= in1[2];
    end
 end
 assign n_1470 = cadence_register_n_1470;
reg cadence_register_n_1471;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1471 <= n_1470;
    end
 end
 assign n_1471 = cadence_register_n_1471;
reg cadence_register_n_1472;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1472 <= in2[18];
    end
 end
 assign n_1472 = cadence_register_n_1472;
reg cadence_register_n_1473;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1473 <= n_1472;
    end
 end
 assign n_1473 = cadence_register_n_1473;
reg cadence_register_n_1474;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1474 <= n_1294;
    end
 end
 assign n_1474 = cadence_register_n_1474;
reg cadence_register_out1_27;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_27 <= n_1474;
    end
 end
 assign out1[27] = cadence_register_out1_27;
reg cadence_register_n_1476;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1476 <= in1_65_2_;
    end
 end
 assign n_1476 = cadence_register_n_1476;
reg cadence_register_n_1477;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1477 <= in2[2];
    end
 end
 assign n_1477 = cadence_register_n_1477;
reg cadence_register_n_1478;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1478 <= n_1477;
    end
 end
 assign n_1478 = cadence_register_n_1478;
reg cadence_register_n_1479;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1479 <= in2[8];
    end
 end
 assign n_1479 = cadence_register_n_1479;
reg cadence_register_n_1480;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1480 <= n_1479;
    end
 end
 assign n_1480 = cadence_register_n_1480;
reg cadence_register_n_1481;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1481 <= in1_65_11_;
    end
 end
 assign n_1481 = cadence_register_n_1481;
reg cadence_register_n_1482;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1482 <= n_1288;
    end
 end
 assign n_1482 = cadence_register_n_1482;
reg cadence_register_out1_33;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_33 <= n_1482;
    end
 end
 assign out1[33] = cadence_register_out1_33;
reg cadence_register_n_1484;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1484 <= in1_43_24_;
    end
 end
 assign n_1484 = cadence_register_n_1484;
reg cadence_register_n_1485;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1485 <= n_1484;
    end
 end
 assign n_1485 = cadence_register_n_1485;
reg cadence_register_n_1486;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1486 <= in1_49_24_;
    end
 end
 assign n_1486 = cadence_register_n_1486;
reg cadence_register_n_1487;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1487 <= n_1486;
    end
 end
 assign n_1487 = cadence_register_n_1487;
reg cadence_register_n_1488;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1488 <= n_1290;
    end
 end
 assign n_1488 = cadence_register_n_1488;
reg cadence_register_out1_31;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_31 <= n_1488;
    end
 end
 assign out1[31] = cadence_register_out1_31;
reg cadence_register_n_1490;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1490 <= in1_65_14_;
    end
 end
 assign n_1490 = cadence_register_n_1490;
reg cadence_register_n_1491;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1491 <= in1_58_24_;
    end
 end
 assign n_1491 = cadence_register_n_1491;
reg cadence_register_n_1492;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1492 <= n_1491;
    end
 end
 assign n_1492 = cadence_register_n_1492;
reg cadence_register_n_1493;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1493 <= in1_61_24_;
    end
 end
 assign n_1493 = cadence_register_n_1493;
reg cadence_register_n_1494;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1494 <= n_1493;
    end
 end
 assign n_1494 = cadence_register_n_1494;
reg cadence_register_n_1495;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1495 <= in2[15];
    end
 end
 assign n_1495 = cadence_register_n_1495;
reg cadence_register_n_1496;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1496 <= n_1495;
    end
 end
 assign n_1496 = cadence_register_n_1496;
reg cadence_register_n_1497;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1497 <= in1_64_15_;
    end
 end
 assign n_1497 = cadence_register_n_1497;
reg cadence_register_n_1498;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1498 <= in1_64_18_;
    end
 end
 assign n_1498 = cadence_register_n_1498;
reg cadence_register_n_1499;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1499 <= in1_65_16_;
    end
 end
 assign n_1499 = cadence_register_n_1499;
reg cadence_register_n_1500;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1500 <= in1_64_17_;
    end
 end
 assign n_1500 = cadence_register_n_1500;
reg cadence_register_n_1501;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1501 <= n_738;
    end
 end
 assign n_1501 = cadence_register_n_1501;
reg cadence_register_n_1502;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1502 <= n_1291;
    end
 end
 assign n_1502 = cadence_register_n_1502;
reg cadence_register_out1_30;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_30 <= n_1502;
    end
 end
 assign out1[30] = cadence_register_out1_30;
reg cadence_register_n_1504;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1504 <= in1_65_9_;
    end
 end
 assign n_1504 = cadence_register_n_1504;
reg cadence_register_n_1505;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1505 <= in1_65_8_;
    end
 end
 assign n_1505 = cadence_register_n_1505;
reg cadence_register_n_1506;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1506 <= in1_65_7_;
    end
 end
 assign n_1506 = cadence_register_n_1506;
reg cadence_register_n_1507;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1507 <= in1_65_6_;
    end
 end
 assign n_1507 = cadence_register_n_1507;
reg cadence_register_n_1508;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1508 <= in1_65_5_;
    end
 end
 assign n_1508 = cadence_register_n_1508;
reg cadence_register_n_1509;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1509 <= in1[10];
    end
 end
 assign n_1509 = cadence_register_n_1509;
reg cadence_register_n_1510;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1510 <= n_1509;
    end
 end
 assign n_1510 = cadence_register_n_1510;
reg cadence_register_n_1511;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1511 <= n_1285;
    end
 end
 assign n_1511 = cadence_register_n_1511;
reg cadence_register_out1_36;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_out1_36 <= n_1511;
    end
 end
 assign out1[36] = cadence_register_out1_36;
reg cadence_register_n_1513;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1513 <= in1_65_10_;
    end
 end
 assign n_1513 = cadence_register_n_1513;
reg cadence_register_n_1514;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1514 <= in1_65_4_;
    end
 end
 assign n_1514 = cadence_register_n_1514;
reg cadence_register_n_1515;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1515 <= in1_65_3_;
    end
 end
 assign n_1515 = cadence_register_n_1515;
reg cadence_register_n_1516;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1516 <= in1_65_13_;
    end
 end
 assign n_1516 = cadence_register_n_1516;
reg cadence_register_n_1517;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1517 <= n_748;
    end
 end
 assign n_1517 = cadence_register_n_1517;
reg cadence_register_n_1518;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1518 <= sub_634_2_n_168;
    end
 end
 assign n_1518 = cadence_register_n_1518;
reg cadence_register_n_1519;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1519 <= n_778;
    end
 end
 assign n_1519 = cadence_register_n_1519;
reg cadence_register_n_1520;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1520 <= sub_634_2_n_23;
    end
 end
 assign n_1520 = cadence_register_n_1520;
reg cadence_register_n_1521;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1521 <= n_737;
    end
 end
 assign n_1521 = cadence_register_n_1521;
reg cadence_register_n_1522;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1522 <= in1[11];
    end
 end
 assign n_1522 = cadence_register_n_1522;
reg cadence_register_n_1523;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1523 <= n_1522;
    end
 end
 assign n_1523 = cadence_register_n_1523;
reg cadence_register_n_1524;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1524 <= n_749;
    end
 end
 assign n_1524 = cadence_register_n_1524;
reg cadence_register_n_1525;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1525 <= n_742;
    end
 end
 assign n_1525 = cadence_register_n_1525;
reg cadence_register_n_1526;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1526 <= in1_65_12_;
    end
 end
 assign n_1526 = cadence_register_n_1526;
reg cadence_register_n_1527;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1527 <= in2[7];
    end
 end
 assign n_1527 = cadence_register_n_1527;
reg cadence_register_n_1528;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1528 <= n_1527;
    end
 end
 assign n_1528 = cadence_register_n_1528;
reg cadence_register_n_1529;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1529 <= in1_65_0_;
    end
 end
 assign n_1529 = cadence_register_n_1529;
reg cadence_register_n_1530;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1530 <= in1[4];
    end
 end
 assign n_1530 = cadence_register_n_1530;
reg cadence_register_n_1531;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1531 <= n_1530;
    end
 end
 assign n_1531 = cadence_register_n_1531;
reg cadence_register_n_1532;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1532 <= in1[18];
    end
 end
 assign n_1532 = cadence_register_n_1532;
reg cadence_register_n_1533;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1533 <= in1_65_1_;
    end
 end
 assign n_1533 = cadence_register_n_1533;
reg cadence_register_n_1534;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1534 <= n_755;
    end
 end
 assign n_1534 = cadence_register_n_1534;
reg cadence_register_n_1535;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1535 <= in2[4];
    end
 end
 assign n_1535 = cadence_register_n_1535;
reg cadence_register_n_1536;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1536 <= n_1535;
    end
 end
 assign n_1536 = cadence_register_n_1536;
reg cadence_register_n_1537;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1537 <= in1[13];
    end
 end
 assign n_1537 = cadence_register_n_1537;
reg cadence_register_n_1538;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1538 <= in1[12];
    end
 end
 assign n_1538 = cadence_register_n_1538;
reg cadence_register_n_1539;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1539 <= n_1538;
    end
 end
 assign n_1539 = cadence_register_n_1539;
reg cadence_register_n_1540;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1540 <= sub_949_2_n_68;
    end
 end
 assign n_1540 = cadence_register_n_1540;
reg cadence_register_n_1541;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1541 <= in1_64_20_;
    end
 end
 assign n_1541 = cadence_register_n_1541;
reg cadence_register_n_1542;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1542 <= in1[23];
    end
 end
 assign n_1542 = cadence_register_n_1542;
reg cadence_register_n_1543;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1543 <= in2[0];
    end
 end
 assign n_1543 = cadence_register_n_1543;
reg cadence_register_n_1544;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1544 <= n_1543;
    end
 end
 assign n_1544 = cadence_register_n_1544;
reg cadence_register_n_1545;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1545 <= sub_655_2_n_82;
    end
 end
 assign n_1545 = cadence_register_n_1545;
reg cadence_register_n_1546;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1546 <= in1[9];
    end
 end
 assign n_1546 = cadence_register_n_1546;
reg cadence_register_n_1547;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1547 <= n_1546;
    end
 end
 assign n_1547 = cadence_register_n_1547;
reg cadence_register_n_1548;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1548 <= in1[14];
    end
 end
 assign n_1548 = cadence_register_n_1548;
reg cadence_register_n_1549;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1549 <= in2[16];
    end
 end
 assign n_1549 = cadence_register_n_1549;
reg cadence_register_n_1550;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1550 <= n_1549;
    end
 end
 assign n_1550 = cadence_register_n_1550;
reg cadence_register_n_1551;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1551 <= in2[10];
    end
 end
 assign n_1551 = cadence_register_n_1551;
reg cadence_register_n_1552;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1552 <= n_1551;
    end
 end
 assign n_1552 = cadence_register_n_1552;
reg cadence_register_n_1553;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1553 <= in1[3];
    end
 end
 assign n_1553 = cadence_register_n_1553;
reg cadence_register_n_1554;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1554 <= n_1553;
    end
 end
 assign n_1554 = cadence_register_n_1554;
reg cadence_register_n_1555;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1555 <= in2[11];
    end
 end
 assign n_1555 = cadence_register_n_1555;
reg cadence_register_n_1556;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1556 <= n_1555;
    end
 end
 assign n_1556 = cadence_register_n_1556;
reg cadence_register_n_1557;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1557 <= in1[17];
    end
 end
 assign n_1557 = cadence_register_n_1557;
reg cadence_register_n_1558;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1558 <= in2[19];
    end
 end
 assign n_1558 = cadence_register_n_1558;
reg cadence_register_n_1559;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1559 <= n_1558;
    end
 end
 assign n_1559 = cadence_register_n_1559;
reg cadence_register_n_1560;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1560 <= in1[16];
    end
 end
 assign n_1560 = cadence_register_n_1560;
reg cadence_register_n_1561;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1561 <= in1[20];
    end
 end
 assign n_1561 = cadence_register_n_1561;
reg cadence_register_n_1562;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1562 <= in2[17];
    end
 end
 assign n_1562 = cadence_register_n_1562;
reg cadence_register_n_1563;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1563 <= n_1562;
    end
 end
 assign n_1563 = cadence_register_n_1563;
reg cadence_register_n_1564;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1564 <= in1[15];
    end
 end
 assign n_1564 = cadence_register_n_1564;
reg cadence_register_n_1565;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1565 <= in2[20];
    end
 end
 assign n_1565 = cadence_register_n_1565;
reg cadence_register_n_1566;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1566 <= n_1565;
    end
 end
 assign n_1566 = cadence_register_n_1566;
reg cadence_register_n_1567;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1567 <= in2[6];
    end
 end
 assign n_1567 = cadence_register_n_1567;
reg cadence_register_n_1568;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1568 <= n_1567;
    end
 end
 assign n_1568 = cadence_register_n_1568;
reg cadence_register_n_1569;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1569 <= in2[5];
    end
 end
 assign n_1569 = cadence_register_n_1569;
reg cadence_register_n_1570;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1570 <= n_1569;
    end
 end
 assign n_1570 = cadence_register_n_1570;
reg cadence_register_n_1571;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1571 <= in1_64_19_;
    end
 end
 assign n_1571 = cadence_register_n_1571;
reg cadence_register_n_1572;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1572 <= in1[24];
    end
 end
 assign n_1572 = cadence_register_n_1572;
reg cadence_register_n_1573;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1573 <= in1[5];
    end
 end
 assign n_1573 = cadence_register_n_1573;
reg cadence_register_n_1574;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1574 <= n_1573;
    end
 end
 assign n_1574 = cadence_register_n_1574;
reg cadence_register_n_1575;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1575 <= in1[6];
    end
 end
 assign n_1575 = cadence_register_n_1575;
reg cadence_register_n_1576;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1576 <= n_1575;
    end
 end
 assign n_1576 = cadence_register_n_1576;
reg cadence_register_n_1577;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1577 <= in2[14];
    end
 end
 assign n_1577 = cadence_register_n_1577;
reg cadence_register_n_1578;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1578 <= n_1577;
    end
 end
 assign n_1578 = cadence_register_n_1578;
reg cadence_register_n_1579;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1579 <= in2[3];
    end
 end
 assign n_1579 = cadence_register_n_1579;
reg cadence_register_n_1580;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1580 <= n_1579;
    end
 end
 assign n_1580 = cadence_register_n_1580;
reg cadence_register_n_1581;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1581 <= in2[13];
    end
 end
 assign n_1581 = cadence_register_n_1581;
reg cadence_register_n_1582;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1582 <= n_1581;
    end
 end
 assign n_1582 = cadence_register_n_1582;
reg cadence_register_n_1583;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1583 <= in1[26];
    end
 end
 assign n_1583 = cadence_register_n_1583;
reg cadence_register_n_1584;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1584 <= in1[19];
    end
 end
 assign n_1584 = cadence_register_n_1584;
reg cadence_register_n_1585;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1585 <= in1[22];
    end
 end
 assign n_1585 = cadence_register_n_1585;
reg cadence_register_n_1586;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1586 <= in2[1];
    end
 end
 assign n_1586 = cadence_register_n_1586;
reg cadence_register_n_1587;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1587 <= n_1586;
    end
 end
 assign n_1587 = cadence_register_n_1587;
reg cadence_register_n_1588;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1588 <= in1[21];
    end
 end
 assign n_1588 = cadence_register_n_1588;
reg cadence_register_n_1589;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1589 <= in2[9];
    end
 end
 assign n_1589 = cadence_register_n_1589;
reg cadence_register_n_1590;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1590 <= n_1589;
    end
 end
 assign n_1590 = cadence_register_n_1590;
reg cadence_register_n_1591;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1591 <= in2[22];
    end
 end
 assign n_1591 = cadence_register_n_1591;
reg cadence_register_n_1592;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1592 <= n_1591;
    end
 end
 assign n_1592 = cadence_register_n_1592;
reg cadence_register_n_1593;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1593 <= in2[21];
    end
 end
 assign n_1593 = cadence_register_n_1593;
reg cadence_register_n_1594;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1594 <= n_1593;
    end
 end
 assign n_1594 = cadence_register_n_1594;
reg cadence_register_n_1595;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1595 <= in2[12];
    end
 end
 assign n_1595 = cadence_register_n_1595;
reg cadence_register_n_1596;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1596 <= n_1595;
    end
 end
 assign n_1596 = cadence_register_n_1596;
reg cadence_register_n_1597;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1597 <= in1[7];
    end
 end
 assign n_1597 = cadence_register_n_1597;
reg cadence_register_n_1598;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1598 <= n_1597;
    end
 end
 assign n_1598 = cadence_register_n_1598;
reg cadence_register_n_1599;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_1599 <= in1[25];
    end
 end
 assign n_1599 = cadence_register_n_1599;
 assign asc001_0_0_ = ~in1_145_24_;
 assign in1_38_12_ = ~(n_1249 & n_1242);
 assign in1_38_9_ = ~(n_1253 & n_1240);
 assign in1_38_6_ = ~(n_1255 & n_1236);
 assign in1_38_5_ = ~(n_1252 & n_1234);
 assign in1_38_8_ = ~(n_1248 & n_1237);
 assign in1_38_4_ = ~(n_1250 & n_1233);
 assign in1_38_0_ = ~(n_1256 & n_1254);
 assign in1_38_11_ = ~(n_1251 & n_1235);
 assign in1_38_10_ = ~(n_1246 & n_1241);
 assign in1_38_7_ = ~(n_1244 & n_1231);
 assign in1_38_2_ = ~(n_1257 & n_1239);
 assign in1_38_1_ = ~(n_1245 & n_1238);
 assign in1_38_3_ = ~(n_1247 & n_1232);
 assign n_1257 = ~(n_1243 & in1_37_2_);
 assign n_1256 = ~(n_1243 & in1_37_0_);
 assign n_1255 = ~(n_1243 & in1_37_6_);
 assign n_1254 = ~(in1_37_24_ & {in1[36]});
 assign n_1253 = ~(in1_37_9_ & ~in1_37_24_);
 assign n_1252 = ~(n_1243 & in1_37_5_);
 assign n_1251 = ~(in1_37_11_ & ~in1_37_24_);
 assign n_1250 = ~(n_1243 & in1_37_4_);
 assign n_1249 = ~(in1_37_12_ & ~in1_37_24_);
 assign n_1248 = ~(n_1243 & in1_37_8_);
 assign n_1247 = ~(n_1243 & in1_37_3_);
 assign n_1246 = ~(n_1243 & in1_37_10_);
 assign n_1245 = ~(n_1243 & in1_37_1_);
 assign n_1244 = ~(n_1243 & in1_37_7_);
 assign n_1243 = ~in1_37_24_;
 assign n_1242 = ~(in1_37_24_ & in1_35_11_);
 assign n_1241 = ~(in1_37_24_ & in1_35_9_);
 assign n_1240 = ~(in1_37_24_ & in1_35_8_);
 assign n_1239 = ~(in1_37_24_ & in1_35_1_);
 assign n_1238 = ~(in1_37_24_ & in1_35_0_);
 assign n_1237 = ~(in1_37_24_ & in1_35_7_);
 assign n_1236 = ~(in1_37_24_ & in1_35_5_);
 assign n_1235 = ~(in1_37_24_ & in1_35_10_);
 assign n_1234 = ~(in1_37_24_ & in1_35_4_);
 assign n_1233 = ~(in1_37_24_ & in1_35_3_);
 assign n_1232 = ~(in1_37_24_ & in1_35_2_);
 assign n_1231 = ~(in1_37_24_ & in1_35_6_);
 assign in1_35_11_ = ~(n_1225 & n_1214);
 assign in1_35_8_ = ~(n_1229 & n_1213);
 assign in1_35_5_ = ~(n_1230 & n_1209);
 assign in1_35_4_ = ~(n_1212 & n_1208);
 assign in1_35_7_ = ~(n_1227 & n_1211);
 assign in1_35_3_ = ~(n_1207 & n_1220);
 assign in1_35_2_ = ~(n_1226 & n_1216);
 assign in1_35_10_ = ~(n_1228 & n_1219);
 assign in1_35_9_ = ~(n_1224 & n_1215);
 assign in1_35_6_ = ~(n_1222 & n_1217);
 assign in1_35_1_ = ~(n_1206 & n_1218);
 assign in1_35_0_ = ~(n_1210 & n_1223);
 assign n_1230 = ~(n_1221 & in1_34_5_);
 assign n_1229 = ~(n_1221 & in1_34_8_);
 assign n_1228 = ~(in1_34_10_ & ~in1_34_24_);
 assign n_1227 = ~(in1_34_7_ & ~in1_34_24_);
 assign n_1226 = ~(n_1221 & in1_34_2_);
 assign n_1225 = ~(in1_34_11_ & ~in1_34_24_);
 assign n_1224 = ~(in1_34_9_ & ~in1_34_24_);
 assign n_1223 = ~(in1_34_24_ & {in1[37]});
 assign n_1222 = ~(n_1221 & in1_34_6_);
 assign n_1221 = ~in1_34_24_;
 assign n_1220 = ~(in1_34_24_ & in1_32_2_);
 assign n_1219 = ~(in1_34_24_ & in1_32_9_);
 assign n_1218 = ~(in1_34_24_ & in1_32_0_);
 assign n_1217 = ~(in1_34_24_ & in1_32_5_);
 assign n_1216 = ~(in1_34_24_ & in1_32_1_);
 assign n_1215 = ~(in1_34_24_ & in1_32_8_);
 assign n_1214 = ~(in1_34_24_ & in1_32_10_);
 assign n_1213 = ~(in1_34_24_ & in1_32_7_);
 assign n_1212 = ~(in1_34_4_ & ~in1_34_24_);
 assign n_1211 = ~(in1_34_24_ & in1_32_6_);
 assign n_1210 = ~(in1_34_0_ & ~in1_34_24_);
 assign n_1209 = ~(in1_34_24_ & in1_32_4_);
 assign n_1208 = ~(in1_34_24_ & in1_32_3_);
 assign n_1207 = ~(in1_34_3_ & ~in1_34_24_);
 assign n_1206 = ~(in1_34_1_ & ~in1_34_24_);
 assign in1_41_5_ = ~(n_1176 & (n_1195 | n_1196));
 assign in1_41_10_ = ~(n_1204 & ~(in1_38_9_ & n_1195));
 assign in1_41_7_ = ~(n_1183 & (n_1188 | n_1194));
 assign in1_41_0_ = ~(n_1205 & (n_1195 | n_1199));
 assign in1_41_6_ = ~(n_1178 & (n_1195 | n_1193));
 assign in1_41_9_ = ~(n_1202 & n_1180);
 assign in1_41_13_ = ~(n_1200 & n_1181);
 assign in1_41_1_ = ~(n_1185 & (n_1188 | n_1190));
 assign in1_41_12_ = ~(n_1186 & (n_1188 | n_1192));
 assign in1_41_11_ = ~(n_1201 & n_1184);
 assign in1_41_8_ = ~(n_1203 & ~(in1_38_7_ & n_1188));
 assign in1_41_3_ = ~(n_1177 & (n_1188 | n_1191));
 assign in1_41_2_ = ~(n_1179 & (n_1195 | n_1197));
 assign in1_41_4_ = ~(n_1182 & (n_1188 | n_1189));
 assign n_1205 = ~(n_1188 & {in1[35]});
 assign n_1204 = ~(n_1187 & in1_40_10_);
 assign n_1203 = (n_1195 | n_1198);
 assign n_1202 = ~(n_1187 & in1_40_9_);
 assign n_1201 = ~(in1_40_11_ & ~n_1195);
 assign n_1200 = ~(in1_40_13_ & ~n_1195);
 assign n_1199 = ~in1_40_0_;
 assign n_1198 = ~in1_40_8_;
 assign n_1197 = ~in1_40_2_;
 assign n_1196 = ~in1_40_5_;
 assign n_1188 = ~n_1187;
 assign n_1195 = ~n_1187;
 assign n_1187 = ~in1_40_24_;
 assign n_1194 = ~in1_40_7_;
 assign n_1193 = ~in1_40_6_;
 assign n_1192 = ~in1_40_12_;
 assign n_1191 = ~in1_40_3_;
 assign n_1190 = ~in1_40_1_;
 assign n_1189 = ~in1_40_4_;
 assign n_1186 = ~(n_1188 & in1_38_11_);
 assign n_1185 = ~(in1_40_24_ & in1_38_0_);
 assign n_1184 = ~(n_1195 & in1_38_10_);
 assign n_1183 = ~(n_1188 & in1_38_6_);
 assign n_1182 = ~(n_1195 & in1_38_3_);
 assign n_1181 = ~(n_1188 & in1_38_12_);
 assign n_1180 = ~(n_1195 & in1_38_8_);
 assign n_1179 = ~(n_1195 & in1_38_1_);
 assign n_1178 = ~(n_1188 & in1_38_5_);
 assign n_1177 = ~(n_1195 & in1_38_2_);
 assign n_1176 = ~(n_1195 & in1_38_4_);
 assign in1_32_4_ = ~(n_1172 & n_1173);
 assign in1_32_7_ = ~(n_1168 & n_1152);
 assign in1_32_10_ = ~(n_1165 & n_1174);
 assign in1_32_3_ = ~(n_1148 & n_1171);
 assign in1_32_6_ = ~(n_1151 & n_1175);
 assign in1_32_2_ = ~(n_1166 & ~(in1_29_1_ & in1_31_24_));
 assign in1_32_1_ = ~(n_1164 & n_1153);
 assign in1_32_9_ = ~(n_1167 & n_1150);
 assign in1_32_8_ = ~(n_1163 & ~(in1_29_7_ & in1_31_24_));
 assign in1_32_5_ = ~(n_1149 & n_1162);
 assign in1_32_0_ = ~(n_1169 & n_1170);
 assign n_1175 = ~(in1_31_24_ & ~n_1159);
 assign n_1174 = ~(in1_31_24_ & ~n_1156);
 assign n_1173 = ~(in1_31_24_ & ~n_1155);
 assign n_1172 = (in1_31_24_ | n_1160);
 assign n_1171 = ~(in1_31_24_ & ~n_1161);
 assign n_1170 = ~(in1_31_24_ & {in1[38]});
 assign n_1169 = ~(n_1154 & in1_31_0_);
 assign n_1168 = ~(n_1154 & in1_31_7_);
 assign n_1167 = ~(in1_31_9_ & n_1154);
 assign n_1166 = (in1_31_24_ | n_1158);
 assign n_1165 = ~(n_1154 & in1_31_10_);
 assign n_1164 = ~(n_1154 & in1_31_1_);
 assign n_1163 = ~(in1_31_8_ & ~in1_31_24_);
 assign n_1162 = ~(in1_31_24_ & ~n_1157);
 assign n_1161 = ~in1_29_2_;
 assign n_1160 = ~in1_31_4_;
 assign n_1159 = ~in1_29_5_;
 assign n_1158 = ~in1_31_2_;
 assign n_1157 = ~in1_29_4_;
 assign n_1156 = ~in1_29_9_;
 assign n_1155 = ~in1_29_3_;
 assign n_1154 = ~in1_31_24_;
 assign n_1153 = ~(in1_31_24_ & in1_29_0_);
 assign n_1152 = ~(in1_31_24_ & in1_29_6_);
 assign n_1151 = ~(in1_31_6_ & ~in1_31_24_);
 assign n_1150 = ~(in1_31_24_ & in1_29_8_);
 assign n_1149 = ~(in1_31_5_ & ~in1_31_24_);
 assign n_1148 = ~(in1_31_3_ & ~in1_31_24_);
 assign in1_44_10_ = ~(n_1142 & ~(in1_41_9_ & in1_43_24_));
 assign in1_44_11_ = ~(n_1146 & n_1126);
 assign in1_44_8_ = ~(n_1147 & ~(in1_41_7_ & in1_43_24_));
 assign in1_44_1_ = ~(n_1131 & n_1122);
 assign in1_44_7_ = ~(n_1125 & n_1133);
 assign in1_44_0_ = ~(n_1119 & ~(in1_43_24_ & {in1[34]}));
 assign in1_44_14_ = ~(n_1143 & n_1132);
 assign in1_44_9_ = ~(n_1128 & n_1121);
 assign in1_44_5_ = ~(n_1124 & n_1123);
 assign in1_44_13_ = ~(n_1145 & n_1127);
 assign in1_44_12_ = ~(n_1141 & n_1135);
 assign in1_44_6_ = ~(n_1144 & ~(in1_41_5_ & in1_43_24_));
 assign in1_44_4_ = ~(n_1129 & n_1130);
 assign in1_44_3_ = ~(n_1118 & n_1120);
 assign in1_44_2_ = ~(n_1134 & n_1136);
 assign n_1147 = (in1_43_24_ | n_1140);
 assign n_1146 = ~(n_1137 & in1_43_11_);
 assign n_1145 = ~(in1_43_13_ & ~in1_43_24_);
 assign n_1144 = (in1_43_24_ | n_1139);
 assign n_1143 = ~(in1_43_14_ & ~in1_43_24_);
 assign n_1142 = (in1_43_24_ | n_1138);
 assign n_1141 = ~(n_1137 & in1_43_12_);
 assign n_1140 = ~in1_43_8_;
 assign n_1139 = ~in1_43_6_;
 assign n_1138 = ~in1_43_10_;
 assign n_1137 = ~in1_43_24_;
 assign n_1136 = ~(in1_43_24_ & in1_41_1_);
 assign n_1135 = ~(in1_43_24_ & in1_41_11_);
 assign n_1134 = ~(in1_43_2_ & ~in1_43_24_);
 assign n_1133 = ~(in1_43_24_ & in1_41_6_);
 assign n_1132 = ~(in1_43_24_ & in1_41_13_);
 assign n_1131 = ~(in1_43_1_ & ~in1_43_24_);
 assign n_1130 = ~(in1_43_24_ & in1_41_3_);
 assign n_1129 = ~(in1_43_4_ & ~in1_43_24_);
 assign n_1128 = ~(in1_43_9_ & ~in1_43_24_);
 assign n_1127 = ~(in1_43_24_ & in1_41_12_);
 assign n_1126 = ~(in1_43_24_ & in1_41_10_);
 assign n_1125 = ~(in1_43_7_ & ~in1_43_24_);
 assign n_1124 = ~(in1_43_5_ & ~in1_43_24_);
 assign n_1123 = ~(in1_43_24_ & in1_41_4_);
 assign n_1122 = ~(in1_43_24_ & in1_41_0_);
 assign n_1121 = ~(in1_43_24_ & in1_41_8_);
 assign n_1120 = ~(in1_43_24_ & in1_41_2_);
 assign n_1119 = ~(in1_43_0_ & ~in1_43_24_);
 assign n_1118 = ~(in1_43_3_ & ~in1_43_24_);
 assign in1_29_3_ = ~(n_1116 & n_1104);
 assign in1_29_6_ = ~(n_1117 & n_1098);
 assign in1_29_9_ = ~(n_1113 & n_1099);
 assign in1_29_2_ = ~(n_1115 & n_1102);
 assign in1_29_5_ = ~(n_1112 & n_1103);
 assign in1_29_8_ = ~(n_1114 & n_1096);
 assign in1_29_0_ = ~(n_1110 & n_1111);
 assign in1_29_1_ = ~(n_1100 & (in1_28_24_ | n_1107));
 assign in1_29_7_ = ~(n_1109 & n_1097);
 assign in1_29_4_ = ~(n_1108 & n_1101);
 assign n_1117 = ~(n_1105 & in1_28_6_);
 assign n_1116 = ~(n_1105 & in1_28_3_);
 assign n_1115 = ~(n_1105 & in1_28_2_);
 assign n_1114 = ~(n_1105 & in1_28_8_);
 assign n_1113 = ~(in1_28_9_ & ~in1_28_24_);
 assign n_1112 = ~(n_1105 & in1_28_5_);
 assign n_1111 = ~(in1_28_24_ & {in1[39]});
 assign n_1110 = ~(n_1105 & in1_28_0_);
 assign n_1109 = ~(n_1105 & in1_28_7_);
 assign n_1108 = (in1_28_24_ | n_1106);
 assign n_1107 = ~in1_28_1_;
 assign n_1106 = ~in1_28_4_;
 assign n_1105 = ~in1_28_24_;
 assign n_1104 = ~(in1_28_24_ & in1_26_2_);
 assign n_1103 = ~(in1_28_24_ & in1_26_4_);
 assign n_1102 = ~(in1_28_24_ & in1_26_1_);
 assign n_1101 = ~(in1_28_24_ & in1_26_3_);
 assign n_1100 = ~(in1_28_24_ & in1_26_0_);
 assign n_1099 = ~(in1_28_24_ & in1_26_8_);
 assign n_1098 = ~(in1_28_24_ & in1_26_5_);
 assign n_1097 = ~(in1_28_24_ & in1_26_6_);
 assign n_1096 = ~(in1_28_24_ & in1_26_7_);
 assign in1_47_8_ = ~(n_1086 & ~(in1_44_7_ & in1_46_24_));
 assign in1_47_12_ = ~(n_1091 & ~(in1_44_11_ & in1_46_24_));
 assign in1_47_9_ = ~(n_1095 & ~(in1_44_8_ & in1_46_24_));
 assign in1_47_2_ = ~(n_1094 & n_1072);
 assign in1_47_15_ = ~(n_1087 & n_1073);
 assign in1_47_1_ = ~(n_1093 & ~(in1_44_0_ & in1_46_24_));
 assign in1_47_0_ = ~(n_1070 & ~(in1_46_24_ & {in1[33]}));
 assign in1_47_11_ = ~(n_1090 & n_1069);
 assign in1_47_10_ = ~(n_1083 & ~(in1_44_9_ & in1_46_24_));
 assign in1_47_6_ = ~(n_1085 & ~(in1_44_5_ & in1_46_24_));
 assign in1_47_14_ = ~(n_1089 & n_1071);
 assign in1_47_13_ = ~(n_1084 & n_1075);
 assign in1_47_7_ = ~(n_1088 & ~(in1_44_6_ & in1_46_24_));
 assign in1_47_5_ = ~(n_1092 & ~(in1_44_4_ & in1_46_24_));
 assign in1_47_4_ = ~(n_1068 & ~(in1_44_3_ & in1_46_24_));
 assign in1_47_3_ = ~(n_1074 & ~(in1_44_2_ & in1_46_24_));
 assign n_1095 = ~(in1_46_9_ & ~in1_46_24_);
 assign n_1094 = (in1_46_24_ | n_1081);
 assign n_1093 = (in1_46_24_ | n_1080);
 assign n_1092 = (in1_46_24_ | n_1078);
 assign n_1091 = ~(in1_46_12_ & ~in1_46_24_);
 assign n_1090 = ~(n_1076 & in1_46_11_);
 assign n_1089 = ~(in1_46_14_ & ~in1_46_24_);
 assign n_1088 = ~(n_1076 & in1_46_7_);
 assign n_1087 = ~(in1_46_15_ & ~in1_46_24_);
 assign n_1086 = (in1_46_24_ | n_1082);
 assign n_1085 = (in1_46_24_ | n_1079);
 assign n_1084 = ~(in1_46_13_ & ~in1_46_24_);
 assign n_1083 = (in1_46_24_ | n_1077);
 assign n_1082 = ~in1_46_8_;
 assign n_1081 = ~in1_46_2_;
 assign n_1080 = ~in1_46_1_;
 assign n_1079 = ~in1_46_6_;
 assign n_1078 = ~in1_46_5_;
 assign n_1077 = ~in1_46_10_;
 assign n_1076 = ~in1_46_24_;
 assign n_1075 = ~(in1_46_24_ & in1_44_12_);
 assign n_1074 = ~(in1_46_3_ & ~in1_46_24_);
 assign n_1073 = ~(in1_46_24_ & in1_44_14_);
 assign n_1072 = ~(in1_46_24_ & in1_44_1_);
 assign n_1071 = ~(in1_46_24_ & in1_44_13_);
 assign n_1070 = ~(in1_46_0_ & ~in1_46_24_);
 assign n_1069 = ~(in1_46_24_ & in1_44_10_);
 assign n_1068 = ~(in1_46_4_ & ~in1_46_24_);
 assign in1_26_2_ = ~(n_1067 & n_1049);
 assign in1_26_5_ = ~(n_1065 & n_1056);
 assign in1_26_8_ = ~(n_1062 & n_1052);
 assign in1_26_1_ = ~(n_1059 & n_1055);
 assign in1_26_7_ = ~(n_1063 & n_1051);
 assign in1_26_0_ = ~(n_1061 & n_1066);
 assign in1_26_4_ = ~(n_1054 & (in1_25_24_ | n_1058));
 assign in1_26_6_ = ~(n_1060 & n_1050);
 assign in1_26_3_ = ~(n_1064 & n_1053);
 assign n_1067 = ~(n_1057 & in1_25_2_);
 assign n_1066 = ~(in1_25_24_ & {in1[40]});
 assign n_1065 = ~(n_1057 & in1_25_5_);
 assign n_1064 = ~(n_1057 & in1_25_3_);
 assign n_1063 = ~(in1_25_7_ & ~in1_25_24_);
 assign n_1062 = ~(in1_25_8_ & ~in1_25_24_);
 assign n_1061 = ~(n_1057 & in1_25_0_);
 assign n_1060 = ~(n_1057 & in1_25_6_);
 assign n_1059 = ~(n_1057 & in1_25_1_);
 assign n_1058 = ~in1_25_4_;
 assign n_1057 = ~in1_25_24_;
 assign n_1056 = ~(in1_25_24_ & in1_23_4_);
 assign n_1055 = ~(in1_25_24_ & in1_23_0_);
 assign n_1054 = ~(in1_25_24_ & in1_23_3_);
 assign n_1053 = ~(in1_25_24_ & in1_23_2_);
 assign n_1052 = ~(in1_25_24_ & in1_23_7_);
 assign n_1051 = ~(in1_25_24_ & in1_23_6_);
 assign n_1050 = ~(in1_25_24_ & in1_23_5_);
 assign n_1049 = ~(in1_25_24_ & in1_23_1_);
 assign in1_50_9_ = ~(n_1046 & n_1021);
 assign in1_50_13_ = ~(n_1043 & n_1022);
 assign in1_50_10_ = ~(n_1047 & n_1030);
 assign in1_50_3_ = ~(n_1028 & n_1029);
 assign in1_50_16_ = ~(n_1039 & n_1020);
 assign in1_50_2_ = ~(n_1026 & n_1027);
 assign in1_50_1_ = ~(n_1048 & ~(in1_47_0_ & in1_49_24_));
 assign in1_50_12_ = ~(n_1044 & n_1018);
 assign in1_50_4_ = ~(n_1017 & ~(in1_47_3_ & in1_49_24_));
 assign in1_50_0_ = ~(n_1041 & n_1045);
 assign in1_50_7_ = ~(n_1016 & (in1_49_24_ | n_1034));
 assign in1_50_15_ = ~(n_1042 & n_1025);
 assign in1_50_14_ = ~(n_1037 & n_1019);
 assign in1_50_11_ = ~(n_1036 & n_1023);
 assign in1_50_6_ = ~(n_1038 & n_1024);
 assign in1_50_5_ = ~(n_1015 & (in1_49_24_ | n_1032));
 assign in1_50_8_ = ~(n_1040 & ~(in1_47_7_ & in1_49_24_));
 assign n_1048 = (in1_49_24_ | n_1033);
 assign n_1047 = ~(n_1031 & in1_49_10_);
 assign n_1046 = ~(n_1031 & in1_49_9_);
 assign n_1045 = ~(in1_49_24_ & {in1[32]});
 assign n_1044 = ~(n_1031 & in1_49_12_);
 assign n_1043 = ~(in1_49_13_ & ~in1_49_24_);
 assign n_1042 = ~(in1_49_15_ & ~in1_49_24_);
 assign n_1041 = ~(n_1031 & in1_49_0_);
 assign n_1040 = (in1_49_24_ | n_1035);
 assign n_1039 = ~(n_1031 & in1_49_16_);
 assign n_1038 = ~(n_1031 & in1_49_6_);
 assign n_1037 = ~(in1_49_14_ & ~in1_49_24_);
 assign n_1036 = ~(in1_49_11_ & ~in1_49_24_);
 assign n_1035 = ~in1_49_8_;
 assign n_1034 = ~in1_49_7_;
 assign n_1033 = ~in1_49_1_;
 assign n_1032 = ~in1_49_5_;
 assign n_1031 = ~in1_49_24_;
 assign n_1030 = ~(in1_49_24_ & in1_47_9_);
 assign n_1029 = ~(in1_49_24_ & in1_47_2_);
 assign n_1028 = ~(in1_49_3_ & ~in1_49_24_);
 assign n_1027 = ~(in1_49_24_ & in1_47_1_);
 assign n_1026 = ~(in1_49_2_ & ~in1_49_24_);
 assign n_1025 = ~(in1_49_24_ & in1_47_14_);
 assign n_1024 = ~(in1_49_24_ & in1_47_5_);
 assign n_1023 = ~(in1_49_24_ & in1_47_10_);
 assign n_1022 = ~(in1_49_24_ & in1_47_12_);
 assign n_1021 = ~(in1_49_24_ & in1_47_8_);
 assign n_1020 = ~(in1_49_24_ & in1_47_15_);
 assign n_1019 = ~(in1_49_24_ & in1_47_13_);
 assign n_1018 = ~(in1_49_24_ & in1_47_11_);
 assign n_1017 = ~(in1_49_4_ & ~in1_49_24_);
 assign n_1016 = ~(in1_49_24_ & in1_47_6_);
 assign n_1015 = ~(in1_49_24_ & in1_47_4_);
 assign in1_23_1_ = ~(n_1014 & ~(in1_20_0_ & in1_22_24_));
 assign in1_23_4_ = ~(n_999 & ~n_1008);
 assign in1_23_7_ = ~(n_1011 & n_1001);
 assign in1_23_0_ = ~(n_1013 & (n_1004 | n_1007));
 assign in1_23_5_ = ~(n_1009 & n_1002);
 assign in1_23_6_ = ~(n_1012 & n_1000);
 assign in1_23_3_ = ~(n_1010 & ~(in1_20_2_ & in1_22_24_));
 assign in1_23_2_ = ~(n_998 & n_997);
 assign n_1014 = (in1_22_24_ | n_1006);
 assign n_1013 = ~(in1_22_24_ & {in1[41]});
 assign n_1012 = ~(in1_22_6_ & ~in1_22_24_);
 assign n_1011 = ~(in1_22_7_ & ~n_1004);
 assign n_1010 = (in1_22_24_ | n_1005);
 assign n_1009 = ~(n_1003 & in1_22_5_);
 assign n_1008 = ~(in1_22_24_ | ~in1_22_4_);
 assign n_1007 = ~in1_22_0_;
 assign n_1006 = ~in1_22_1_;
 assign n_1005 = ~in1_22_3_;
 assign n_1004 = ~n_1003;
 assign n_1003 = ~in1_22_24_;
 assign n_1002 = ~(n_1004 & in1_20_4_);
 assign n_1001 = ~(n_1004 & in1_20_6_);
 assign n_1000 = ~(n_1004 & in1_20_5_);
 assign n_999 = ~(n_1004 & in1_20_3_);
 assign n_998 = ~(in1_22_2_ & ~in1_22_24_);
 assign n_997 = ~(n_1004 & in1_20_1_);
 assign in1_53_9_ = ~(n_962 & n_972);
 assign in1_53_14_ = ~(n_992 & n_976);
 assign in1_53_11_ = ~(n_996 & n_977);
 assign in1_53_4_ = ~(n_995 & n_971);
 assign in1_53_10_ = ~(n_993 & n_978);
 assign in1_53_3_ = ~(n_980 & ~n_994);
 assign in1_53_2_ = ~(n_973 & n_974);
 assign in1_53_13_ = ~(n_989 & n_975);
 assign in1_53_17_ = ~(n_990 & n_982);
 assign in1_53_5_ = ~(n_963 & n_960);
 assign in1_53_0_ = ~(n_981 & n_991);
 assign in1_53_8_ = ~(n_961 & n_966);
 assign in1_53_16_ = ~(n_970 & (in1_52_24_ | n_986));
 assign in1_53_15_ = ~(n_988 & n_983);
 assign in1_53_12_ = ~(n_987 & n_964);
 assign in1_53_7_ = ~(n_967 & ~(n_985 & in1_52_7_));
 assign in1_53_6_ = ~(n_965 & n_979);
 assign in1_53_1_ = ~(n_968 & ~n_969);
 assign n_996 = ~(n_985 & in1_52_11_);
 assign n_995 = ~(n_985 & in1_52_4_);
 assign n_994 = ~(in1_52_24_ | ~in1_52_3_);
 assign n_993 = ~(n_985 & in1_52_10_);
 assign n_992 = ~(n_985 & in1_52_14_);
 assign n_991 = ~(in1_52_24_ & {in1[31]});
 assign n_990 = ~(in1_52_17_ & ~in1_52_24_);
 assign n_989 = ~(n_985 & in1_52_13_);
 assign n_988 = ~(in1_52_15_ & ~in1_52_24_);
 assign n_987 = (in1_52_24_ | n_984);
 assign n_986 = ~in1_52_16_;
 assign n_985 = ~in1_52_24_;
 assign n_984 = ~in1_52_12_;
 assign n_983 = ~(in1_52_24_ & in1_50_14_);
 assign n_982 = ~(in1_52_24_ & in1_50_16_);
 assign n_981 = ~(in1_52_0_ & ~in1_52_24_);
 assign n_980 = ~(in1_52_24_ & in1_50_2_);
 assign n_979 = ~(in1_52_24_ & in1_50_5_);
 assign n_978 = ~(in1_52_24_ & in1_50_9_);
 assign n_977 = ~(in1_52_24_ & in1_50_10_);
 assign n_976 = ~(in1_52_24_ & in1_50_13_);
 assign n_975 = ~(in1_52_24_ & in1_50_12_);
 assign n_974 = ~(in1_52_24_ & in1_50_1_);
 assign n_973 = ~(in1_52_2_ & ~in1_52_24_);
 assign n_972 = ~(in1_52_24_ & in1_50_8_);
 assign n_971 = ~(in1_52_24_ & in1_50_3_);
 assign n_970 = ~(in1_52_24_ & in1_50_15_);
 assign n_969 = ~(in1_52_24_ | ~in1_52_1_);
 assign n_968 = ~(in1_52_24_ & in1_50_0_);
 assign n_967 = ~(in1_52_24_ & in1_50_6_);
 assign n_966 = ~(in1_52_24_ & in1_50_7_);
 assign n_965 = ~(in1_52_6_ & ~in1_52_24_);
 assign n_964 = ~(in1_52_24_ & in1_50_11_);
 assign n_963 = ~(in1_52_5_ & ~in1_52_24_);
 assign n_962 = ~(in1_52_9_ & ~in1_52_24_);
 assign n_961 = ~(in1_52_8_ & ~in1_52_24_);
 assign n_960 = ~(in1_52_24_ & in1_50_4_);
 assign in1_20_6_ = ~(n_956 & n_952);
 assign in1_20_3_ = ~(n_951 & ~(in1_17_2_ & in1_19_24_));
 assign in1_20_0_ = ~(n_958 & n_959);
 assign in1_20_4_ = ~(n_946 & n_948);
 assign in1_20_5_ = ~(n_957 & n_947);
 assign in1_20_2_ = ~(n_955 & ~(in1_17_1_ & in1_19_24_));
 assign in1_20_1_ = ~(n_950 & n_949);
 assign n_959 = ~(in1_19_24_ & {in1[42]});
 assign n_958 = (in1_19_24_ | n_954);
 assign n_957 = ~(in1_19_5_ & ~in1_19_24_);
 assign n_956 = ~(in1_19_6_ & ~in1_19_24_);
 assign n_955 = (in1_19_24_ | n_953);
 assign n_954 = ~in1_19_0_;
 assign n_953 = ~in1_19_2_;
 assign n_952 = ~(in1_19_24_ & in1_17_5_);
 assign n_951 = ~(in1_19_3_ & ~in1_19_24_);
 assign n_950 = ~(in1_19_1_ & ~in1_19_24_);
 assign n_949 = ~(in1_19_24_ & in1_17_0_);
 assign n_948 = ~(in1_19_24_ & in1_17_3_);
 assign n_947 = ~(in1_19_24_ & in1_17_4_);
 assign n_946 = ~(in1_19_4_ & ~in1_19_24_);
 assign in1_56_10_ = ~(n_941 & n_913);
 assign in1_56_15_ = ~(n_938 & n_925);
 assign in1_56_12_ = ~(n_916 & n_910);
 assign in1_56_5_ = ~(n_945 & n_917);
 assign in1_56_11_ = ~(n_928 & n_914);
 assign in1_56_4_ = ~(n_926 & n_909);
 assign in1_56_3_ = ~(n_921 & n_924);
 assign in1_56_14_ = ~(n_937 & n_907);
 assign in1_56_18_ = ~(n_939 & n_927);
 assign in1_56_2_ = ~(n_905 & n_920);
 assign in1_56_1_ = ~(n_904 & n_912);
 assign in1_56_9_ = ~(n_936 & n_911);
 assign in1_56_0_ = ~(n_943 & n_944);
 assign in1_56_17_ = ~(n_942 & n_915);
 assign in1_56_16_ = ~(n_935 & n_919);
 assign in1_56_13_ = ~(n_922 & ~(n_932 & in1_55_13_));
 assign in1_56_8_ = ~(n_940 & n_906);
 assign in1_56_7_ = ~(n_918 & ~n_934);
 assign in1_56_6_ = ~(n_923 & n_908);
 assign n_945 = ~(n_932 & in1_55_5_);
 assign n_944 = ~(in1_55_24_ & {in1[30]});
 assign n_943 = ~(n_932 & in1_55_0_);
 assign n_942 = ~(n_932 & in1_55_17_);
 assign n_941 = (in1_55_24_ | n_933);
 assign n_940 = (in1_55_24_ | n_929);
 assign n_939 = ~(n_932 & in1_55_18_);
 assign n_938 = ~(in1_55_15_ & ~in1_55_24_);
 assign n_937 = ~(n_932 & in1_55_14_);
 assign n_936 = (in1_55_24_ | n_930);
 assign n_935 = (in1_55_24_ | n_931);
 assign n_934 = ~(in1_55_24_ | ~in1_55_7_);
 assign n_933 = ~in1_55_10_;
 assign n_932 = ~in1_55_24_;
 assign n_931 = ~in1_55_16_;
 assign n_930 = ~in1_55_9_;
 assign n_929 = ~in1_55_8_;
 assign n_928 = ~(in1_55_11_ & ~in1_55_24_);
 assign n_927 = ~(in1_55_24_ & in1_53_17_);
 assign n_926 = ~(in1_55_4_ & ~in1_55_24_);
 assign n_925 = ~(in1_55_24_ & in1_53_14_);
 assign n_924 = ~(in1_55_24_ & in1_53_2_);
 assign n_923 = ~(in1_55_6_ & ~in1_55_24_);
 assign n_922 = ~(in1_55_24_ & in1_53_12_);
 assign n_921 = ~(in1_55_3_ & ~in1_55_24_);
 assign n_920 = ~(in1_55_24_ & in1_53_1_);
 assign n_919 = ~(in1_55_24_ & in1_53_15_);
 assign n_918 = ~(in1_55_24_ & in1_53_6_);
 assign n_917 = ~(in1_55_24_ & in1_53_4_);
 assign n_916 = ~(in1_55_12_ & ~in1_55_24_);
 assign n_915 = ~(in1_55_24_ & in1_53_16_);
 assign n_914 = ~(in1_55_24_ & in1_53_10_);
 assign n_913 = ~(in1_55_24_ & in1_53_9_);
 assign n_912 = ~(in1_55_24_ & in1_53_0_);
 assign n_911 = ~(in1_55_24_ & in1_53_8_);
 assign n_910 = ~(in1_55_24_ & in1_53_11_);
 assign n_909 = ~(in1_55_24_ & in1_53_3_);
 assign n_908 = ~(in1_55_24_ & in1_53_5_);
 assign n_907 = ~(in1_55_24_ & in1_53_13_);
 assign n_906 = ~(in1_55_24_ & in1_53_7_);
 assign n_905 = ~(in1_55_2_ & ~in1_55_24_);
 assign n_904 = ~(in1_55_1_ & ~in1_55_24_);
 assign in1_17_5_ = ~(n_891 & (n_897 | n_900));
 assign in1_17_2_ = ~(n_902 & ~(in1_14_1_ & in1_16_24_));
 assign in1_17_1_ = ~(n_893 & (n_897 | n_898));
 assign in1_17_4_ = ~(n_903 & n_895);
 assign in1_17_3_ = ~(n_890 & n_894);
 assign in1_17_0_ = ~(n_892 & n_901);
 assign n_903 = ~(n_896 & in1_16_4_);
 assign n_902 = (in1_16_24_ | n_899);
 assign n_901 = ~(in1_16_24_ & {in1[43]});
 assign n_900 = ~in1_16_5_;
 assign n_899 = ~in1_16_2_;
 assign n_898 = ~in1_16_1_;
 assign n_897 = ~n_896;
 assign n_896 = ~in1_16_24_;
 assign n_895 = ~(in1_16_24_ & in1_14_3_);
 assign n_894 = ~(in1_16_24_ & in1_14_2_);
 assign n_893 = ~(n_897 & in1_14_0_);
 assign n_892 = ~(in1_16_0_ & ~in1_16_24_);
 assign n_891 = ~(n_897 & in1_14_4_);
 assign n_890 = ~(in1_16_3_ & ~in1_16_24_);
 assign in1_59_19_ = ~(n_881 & n_855);
 assign in1_59_16_ = ~(n_884 & n_863);
 assign in1_59_13_ = ~(n_856 & (in1_58_24_ | n_867));
 assign in1_59_6_ = ~(n_888 & ~(in1_56_5_ & in1_58_24_));
 assign in1_59_12_ = ~(n_886 & n_849);
 assign in1_59_5_ = ~(n_887 & n_854);
 assign in1_59_4_ = ~(n_885 & ~(in1_56_3_ & in1_58_24_));
 assign in1_59_15_ = ~(n_880 & n_862);
 assign in1_59_11_ = ~(n_865 & n_860);
 assign in1_59_3_ = ~(n_861 & (in1_58_24_ | n_871));
 assign in1_59_2_ = ~(n_882 & n_851);
 assign in1_59_10_ = ~(n_852 & n_850);
 assign in1_59_1_ = ~(n_847 & (in1_58_24_ | n_875));
 assign in1_59_18_ = ~(n_883 & n_864);
 assign in1_59_17_ = ~(n_878 & n_858);
 assign in1_59_0_ = ~((in1_58_24_ | n_868) & (n_866 | n_873));
 assign in1_59_14_ = ~(n_876 & n_857);
 assign in1_59_9_ = ~(n_879 & n_859);
 assign in1_59_8_ = ~(n_877 & n_848);
 assign in1_59_7_ = ~(n_889 & n_853);
 assign n_889 = ~(n_866 & in1_58_7_);
 assign n_888 = (in1_58_24_ | n_874);
 assign n_887 = ~(n_866 & in1_58_5_);
 assign n_886 = ~(n_866 & in1_58_12_);
 assign n_885 = (in1_58_24_ | n_872);
 assign n_884 = (in1_58_24_ | n_870);
 assign n_883 = ~(in1_58_18_ & ~in1_58_24_);
 assign n_882 = ~(n_866 & in1_58_2_);
 assign n_881 = ~(in1_58_19_ & ~in1_58_24_);
 assign n_880 = ~(n_866 & in1_58_15_);
 assign n_879 = ~(n_866 & in1_58_9_);
 assign n_878 = ~(n_866 & in1_58_17_);
 assign n_877 = (in1_58_24_ | n_869);
 assign n_876 = ~(n_866 & in1_58_14_);
 assign n_875 = ~in1_58_1_;
 assign n_874 = ~in1_58_6_;
 assign n_873 = ~{in1[29]};
 assign n_872 = ~in1_58_4_;
 assign n_871 = ~in1_58_3_;
 assign n_870 = ~in1_58_16_;
 assign n_869 = ~in1_58_8_;
 assign n_868 = ~in1_58_0_;
 assign n_867 = ~in1_58_13_;
 assign n_866 = ~in1_58_24_;
 assign n_865 = ~(in1_58_11_ & ~in1_58_24_);
 assign n_864 = ~(in1_58_24_ & in1_56_17_);
 assign n_863 = ~(in1_58_24_ & in1_56_15_);
 assign n_862 = ~(in1_58_24_ & in1_56_14_);
 assign n_861 = ~(in1_58_24_ & in1_56_2_);
 assign n_860 = ~(in1_58_24_ & in1_56_10_);
 assign n_859 = ~(in1_58_24_ & in1_56_8_);
 assign n_858 = ~(in1_58_24_ & in1_56_16_);
 assign n_857 = ~(in1_58_24_ & in1_56_13_);
 assign n_856 = ~(in1_58_24_ & in1_56_12_);
 assign n_855 = ~(in1_58_24_ & in1_56_18_);
 assign n_854 = ~(in1_58_24_ & in1_56_4_);
 assign n_853 = ~(in1_58_24_ & in1_56_6_);
 assign n_852 = ~(in1_58_10_ & ~in1_58_24_);
 assign n_851 = ~(in1_58_24_ & in1_56_1_);
 assign n_850 = ~(in1_58_24_ & in1_56_9_);
 assign n_849 = ~(in1_58_24_ & in1_56_11_);
 assign n_848 = ~(in1_58_24_ & in1_56_7_);
 assign n_847 = ~(in1_58_24_ & in1_56_0_);
 assign in1_14_4_ = ~(n_844 & n_835);
 assign in1_14_1_ = ~(n_838 & n_840);
 assign in1_14_0_ = ~(n_839 & n_846);
 assign in1_14_3_ = ~(n_845 & n_837);
 assign in1_14_2_ = ~(n_843 & n_836);
 assign n_846 = ~(in1_13_24_ & {in1[44]});
 assign n_845 = ~(n_841 & in1_13_3_);
 assign n_844 = ~(n_841 & in1_13_4_);
 assign n_843 = (in1_13_24_ | n_842);
 assign n_842 = ~in1_13_2_;
 assign n_841 = ~in1_13_24_;
 assign n_840 = ~(in1_13_24_ & in1_11_0_);
 assign n_839 = ~(in1_13_0_ & ~in1_13_24_);
 assign n_838 = ~(in1_13_1_ & ~in1_13_24_);
 assign n_837 = ~(in1_13_24_ & in1_11_2_);
 assign n_836 = ~(in1_13_24_ & in1_11_1_);
 assign n_835 = ~(in1_13_24_ & in1_11_3_);
 assign in1_62_20_ = ~(n_825 & n_791);
 assign in1_62_17_ = ~(n_829 & n_796);
 assign in1_62_14_ = ~(n_832 & n_798);
 assign in1_62_7_ = ~(n_797 & n_800);
 assign in1_62_13_ = ~(n_831 & n_808);
 assign in1_62_6_ = ~(n_790 & n_809);
 assign in1_62_5_ = ~(n_830 & n_795);
 assign in1_62_16_ = ~(n_824 & n_807);
 assign in1_62_12_ = ~(n_811 & ~(n_812 & in1_61_12_));
 assign in1_62_4_ = ~(n_828 & n_806);
 assign in1_62_1_ = ~(n_787 & n_789);
 assign in1_62_11_ = ~(n_821 & n_810);
 assign in1_62_2_ = ~(n_823 & n_794);
 assign in1_62_19_ = ~(n_827 & n_788);
 assign in1_62_18_ = ~(n_819 & n_799);
 assign in1_62_3_ = ~(n_805 & n_803);
 assign in1_62_0_ = ~(n_820 & n_834);
 assign in1_62_15_ = ~(n_826 & n_801);
 assign in1_62_10_ = ~(n_822 & n_802);
 assign in1_62_9_ = ~(n_793 & n_804);
 assign in1_62_8_ = ~(n_833 & n_792);
 assign n_834 = ~(in1_61_24_ & {in1[28]});
 assign n_833 = (n_814 | n_816);
 assign n_832 = ~(n_812 & in1_61_14_);
 assign n_831 = ~(n_812 & in1_61_13_);
 assign n_830 = ~(n_812 & in1_61_5_);
 assign n_829 = ~(n_812 & in1_61_17_);
 assign n_828 = ~(n_812 & in1_61_4_);
 assign n_827 = ~(in1_61_19_ & ~n_813);
 assign n_826 = ~(in1_61_15_ & ~n_813);
 assign n_825 = ~(n_812 & in1_61_20_);
 assign n_824 = (n_813 | n_818);
 assign n_823 = ~(n_815 & in1_61_2_);
 assign n_822 = (n_814 | n_817);
 assign n_821 = ~(n_812 & in1_61_11_);
 assign n_820 = ~(n_815 & in1_61_0_);
 assign n_819 = ~(in1_61_18_ & ~n_813);
 assign n_818 = ~in1_61_16_;
 assign n_817 = ~in1_61_10_;
 assign n_816 = ~in1_61_8_;
 assign n_814 = ~n_815;
 assign n_815 = ~in1_61_24_;
 assign n_813 = ~n_812;
 assign n_812 = ~in1_61_24_;
 assign n_811 = ~(in1_61_24_ & in1_59_11_);
 assign n_810 = ~(n_814 & in1_59_10_);
 assign n_809 = ~(in1_61_24_ & in1_59_5_);
 assign n_808 = ~(n_814 & in1_59_12_);
 assign n_807 = ~(n_813 & in1_59_15_);
 assign n_806 = ~(in1_61_24_ & in1_59_3_);
 assign n_805 = ~(in1_61_3_ & ~in1_61_24_);
 assign n_804 = ~(n_814 & in1_59_8_);
 assign n_803 = ~(n_814 & in1_59_2_);
 assign n_802 = ~(n_814 & in1_59_9_);
 assign n_801 = ~(n_813 & in1_59_14_);
 assign n_800 = ~(n_814 & in1_59_6_);
 assign n_799 = ~(n_813 & in1_59_17_);
 assign n_798 = ~(n_814 & in1_59_13_);
 assign n_797 = ~(in1_61_7_ & ~n_814);
 assign n_796 = ~(n_813 & in1_59_16_);
 assign n_795 = ~(n_814 & in1_59_4_);
 assign n_794 = ~(in1_61_24_ & in1_59_1_);
 assign n_793 = ~(in1_61_9_ & ~in1_61_24_);
 assign n_792 = ~(n_814 & in1_59_7_);
 assign n_791 = ~(n_813 & in1_59_19_);
 assign n_790 = ~(in1_61_6_ & ~in1_61_24_);
 assign n_789 = ~(in1_61_24_ & in1_59_0_);
 assign n_788 = ~(n_813 & in1_59_18_);
 assign n_787 = ~(in1_61_1_ & ~in1_61_24_);
 assign in1_11_3_ = ~(n_785 & (n_786 | in1_10_24_));
 assign in1_11_0_ = ~(n_783 & ~(in1_10_24_ & {in1[45]}));
 assign in1_11_2_ = ~(n_784 & n_782);
 assign in1_11_1_ = ~(n_781 & n_780);
 assign n_786 = ~in1_10_3_;
 assign n_785 = ~(in1_10_24_ & in1_8_2_);
 assign n_784 = ~(in1_10_2_ & ~in1_10_24_);
 assign n_783 = ~(in1_10_0_ & ~in1_10_24_);
 assign n_782 = ~(in1_10_24_ & in1_8_1_);
 assign n_781 = ~(in1_10_1_ & ~in1_10_24_);
 assign n_780 = ~(in1_10_24_ & in1_8_0_);
 assign in1_65_7_ = ~(n_741 & (n_755 | n_754));
 assign in1_65_18_ = ~(n_772 & n_1524);
 assign in1_65_15_ = ~(n_777 & n_1517);
 assign in1_65_8_ = ~(n_776 & n_750);
 assign in1_65_14_ = ~(n_774 & n_732);
 assign in1_65_21_ = ~(n_768 & n_1525);
 assign in1_65_6_ = ~(n_773 & n_735);
 assign in1_65_17_ = ~(n_767 & n_1501);
 assign in1_65_13_ = ~(n_770 & n_739);
 assign in1_65_5_ = ~(n_734 & n_740);
 assign in1_65_4_ = ~(n_769 & n_747);
 assign in1_65_1_ = ~(n_744 & (in1_64_24_ | n_759));
 assign in1_65_3_ = ~(n_745 & (n_755 | n_756));
 assign in1_65_20_ = ~(n_771 & n_1519);
 assign in1_65_19_ = ~(n_762 & n_1521);
 assign in1_65_2_ = ~(n_766 & n_731);
 assign in1_65_12_ = ~(n_765 & ~(in1_62_11_ & n_755));
 assign in1_65_16_ = ~(n_761 & n_733);
 assign in1_65_11_ = ~(n_763 & ~(in1_62_10_ & n_755));
 assign in1_65_0_ = ~(n_775 & n_764);
 assign in1_65_10_ = ~(n_746 & n_736);
 assign in1_65_9_ = ~(n_779 & n_743);
 assign n_779 = ~(n_752 & in1_64_9_);
 assign n_778 = ~(in1_62_19_ & n_755);
 assign n_777 = ~(n_1497 & ~n_1534);
 assign n_776 = (in1_64_24_ | n_760);
 assign n_775 = ~(n_752 & in1_64_0_);
 assign n_774 = ~(in1_64_14_ & ~n_751);
 assign n_773 = (n_751 | n_757);
 assign n_772 = ~(n_1498 & ~n_1534);
 assign n_771 = ~(n_1541 & ~n_1534);
 assign n_770 = ~(in1_64_13_ & ~n_755);
 assign n_769 = (n_751 | n_753);
 assign n_768 = ~(in1_64_21_ & ~n_1534);
 assign n_767 = ~(n_1500 & ~n_1534);
 assign n_766 = ~(n_752 & in1_64_2_);
 assign n_765 = (n_755 | n_758);
 assign n_764 = ~(in1_64_24_ & {in1[27]});
 assign n_763 = ~(n_752 & in1_64_11_);
 assign n_762 = ~(n_1571 & ~n_1534);
 assign n_761 = ~(n_752 & in1_64_16_);
 assign n_760 = ~in1_64_8_;
 assign n_759 = ~in1_64_1_;
 assign n_758 = ~in1_64_12_;
 assign n_757 = ~in1_64_6_;
 assign n_756 = ~in1_64_3_;
 assign n_755 = ~n_752;
 assign n_751 = ~n_752;
 assign n_752 = ~in1_64_24_;
 assign n_754 = ~in1_64_7_;
 assign n_753 = ~in1_64_4_;
 assign n_750 = ~(n_751 & in1_62_7_);
 assign n_749 = ~(n_755 & in1_62_17_);
 assign n_748 = ~(n_755 & in1_62_14_);
 assign n_747 = ~(n_751 & in1_62_3_);
 assign n_746 = ~(in1_64_10_ & ~n_751);
 assign n_745 = ~(n_755 & in1_62_2_);
 assign n_744 = ~(in1_64_24_ & in1_62_0_);
 assign n_743 = ~(n_751 & in1_62_8_);
 assign n_742 = ~(n_755 & in1_62_20_);
 assign n_741 = ~(n_751 & in1_62_6_);
 assign n_740 = ~(n_751 & in1_62_4_);
 assign n_739 = ~(n_755 & in1_62_12_);
 assign n_738 = ~(n_755 & in1_62_16_);
 assign n_737 = ~(n_755 & in1_62_18_);
 assign n_736 = ~(n_751 & in1_62_9_);
 assign n_735 = ~(n_755 & in1_62_5_);
 assign n_734 = ~(in1_64_5_ & ~in1_64_24_);
 assign n_733 = ~(n_755 & in1_62_15_);
 assign n_732 = ~(n_751 & in1_62_13_);
 assign n_731 = ~(in1_64_24_ & in1_62_1_);
 assign in1_8_2_ = ~(n_730 & n_728);
 assign in1_8_1_ = ~(n_727 & n_729);
 assign in1_8_0_ = ~(n_726 & ~(in1_7_24_ & {in1[46]}));
 assign n_730 = ~(in1_7_2_ & ~in1_7_24_);
 assign n_729 = ~(in1_7_24_ & in1_5_0_);
 assign n_728 = ~(in1_7_24_ & in1_5_1_);
 assign n_727 = ~(in1_7_1_ & ~in1_7_24_);
 assign n_726 = ~(in1_7_0_ & ~in1_7_24_);
 assign in1_68_8_ = ~(n_721 & n_694);
 assign in1_68_19_ = ~(n_717 & n_692);
 assign in1_68_16_ = ~(n_724 & n_672);
 assign in1_68_9_ = ~(n_695 & n_677);
 assign in1_68_15_ = ~(n_719 & n_682);
 assign in1_68_22_ = ~(n_713 & n_683);
 assign in1_68_7_ = ~(n_718 & n_691);
 assign in1_68_18_ = ~(n_712 & n_673);
 assign in1_68_14_ = ~(n_715 & n_689);
 assign in1_68_6_ = ~(n_716 & n_722);
 assign in1_68_5_ = ~(n_714 & n_675);
 assign in1_68_17_ = ~(n_679 & ~(n_706 & in1_67_17_));
 assign in1_68_4_ = ~(n_723 & n_688);
 assign in1_68_21_ = ~(n_711 & n_676);
 assign in1_68_20_ = ~(n_709 & n_690);
 assign in1_68_3_ = ~(n_687 & n_685);
 assign in1_68_2_ = ~(n_671 & n_696);
 assign in1_68_13_ = ~(n_686 & ~(n_706 & in1_67_13_));
 assign in1_68_12_ = ~(n_710 & n_693);
 assign in1_68_1_ = ~(n_720 & n_681);
 assign in1_68_11_ = ~(n_680 & n_684);
 assign in1_68_0_ = ~(n_708 & n_725);
 assign in1_68_10_ = ~(n_674 & n_678);
 assign n_725 = ~(in1_67_24_ & n_1583);
 assign n_724 = ~(n_706 & in1_67_16_);
 assign n_723 = (in1_67_24_ | n_701);
 assign n_722 = ~(n_705 & ~n_699);
 assign n_721 = (n_704 | n_700);
 assign n_720 = ~(n_702 & in1_67_1_);
 assign n_719 = ~(n_697 & ~n_703);
 assign n_718 = (n_704 | n_698);
 assign n_717 = ~(in1_67_19_ & ~n_703);
 assign n_716 = ~(n_706 & in1_67_6_);
 assign n_715 = ~(in1_67_14_ & ~n_704);
 assign n_714 = ~(n_706 & in1_67_5_);
 assign n_713 = ~(in1_67_22_ & ~n_703);
 assign n_712 = ~(n_706 & in1_67_18_);
 assign n_711 = ~(in1_67_21_ & ~n_703);
 assign n_710 = (n_704 | n_707);
 assign n_709 = ~(in1_67_20_ & ~n_703);
 assign n_708 = ~(n_706 & in1_67_0_);
 assign n_707 = ~in1_67_12_;
 assign n_705 = ~n_706;
 assign n_703 = ~n_706;
 assign n_704 = ~n_706;
 assign n_706 = ~in1_67_24_;
 assign n_702 = ~in1_67_24_;
 assign n_701 = ~in1_67_4_;
 assign n_700 = ~in1_67_8_;
 assign n_699 = ~n_1508;
 assign n_698 = ~in1_67_7_;
 assign n_697 = in1_67_15_;
 assign n_696 = ~(in1_67_24_ & n_1533);
 assign n_695 = ~(in1_67_9_ & ~n_704);
 assign n_694 = ~(n_704 & n_1506);
 assign n_693 = ~(n_704 & n_1481);
 assign n_692 = ~(n_703 & in1_65_18_);
 assign n_691 = ~(n_704 & n_1507);
 assign n_690 = ~(n_703 & in1_65_19_);
 assign n_689 = ~(n_704 & n_1516);
 assign n_688 = ~(in1_67_24_ & n_1515);
 assign n_687 = ~(in1_67_3_ & ~in1_67_24_);
 assign n_686 = ~(n_704 & n_1526);
 assign n_685 = ~(in1_67_24_ & n_1476);
 assign n_684 = ~(n_704 & n_1513);
 assign n_683 = ~(n_703 & in1_65_21_);
 assign n_682 = ~(n_703 & n_1490);
 assign n_681 = ~(in1_67_24_ & n_1529);
 assign n_680 = ~(in1_67_11_ & ~n_704);
 assign n_679 = ~(n_704 & n_1499);
 assign n_678 = ~(n_704 & n_1504);
 assign n_677 = ~(n_704 & n_1505);
 assign n_676 = ~(n_703 & in1_65_20_);
 assign n_675 = ~(in1_67_24_ & n_1514);
 assign n_674 = ~(in1_67_10_ & ~n_704);
 assign n_673 = ~(n_703 & in1_65_17_);
 assign n_672 = ~(n_704 & in1_65_15_);
 assign n_671 = ~(in1_67_2_ & ~in1_67_24_);
 assign in1_5_1_ = ~(n_665 & n_668);
 assign in1_5_0_ = ~(n_670 & n_669);
 assign n_670 = (in1_4_24_ | n_667);
 assign n_669 = ~(in1_4_24_ & {in1[47]});
 assign n_668 = ~(n_666 & in1_4_1_);
 assign n_667 = ~in1_4_0_;
 assign n_666 = ~in1_4_24_;
 assign n_665 = ~(in1_4_24_ & in1_2_0_);
 assign in1_71_8_ = ~(n_658 & n_624);
 assign in1_71_20_ = ~(n_657 & n_635);
 assign in1_71_17_ = ~(n_661 & ~(in1_68_16_ & in1_70_24_));
 assign in1_71_10_ = ~(n_660 & n_620);
 assign in1_71_16_ = ~(n_659 & n_634);
 assign in1_71_9_ = ~(n_625 & n_616);
 assign in1_71_23_ = ~(n_655 & ~(n_640 & in1_70_23_));
 assign in1_71_19_ = ~(n_653 & n_654);
 assign in1_71_15_ = ~(n_664 & n_615);
 assign in1_71_7_ = ~(n_632 & n_633);
 assign in1_71_6_ = ~(n_630 & n_618);
 assign in1_71_14_ = ~(n_651 & n_628);
 assign in1_71_13_ = ~(n_650 & n_614);
 assign in1_71_22_ = ~(n_656 & n_619);
 assign in1_71_21_ = ~(n_648 & n_631);
 assign in1_71_4_ = ~(n_627 & n_623);
 assign in1_71_3_ = ~(n_626 & (in1_70_24_ | n_637));
 assign in1_71_18_ = ~(n_645 & ~(in1_68_17_ & in1_70_24_));
 assign in1_71_5_ = ~(n_662 & n_617);
 assign in1_71_2_ = ~(n_652 & n_636);
 assign in1_71_12_ = ~(n_647 & n_622);
 assign in1_71_1_ = ~(n_629 & (in1_70_24_ | n_642));
 assign in1_71_0_ = ~(n_646 & n_649);
 assign in1_71_11_ = ~(n_663 & n_621);
 assign n_664 = ~(in1_70_15_ & ~in1_70_24_);
 assign n_663 = (in1_70_24_ | n_641);
 assign n_662 = (in1_70_24_ | n_638);
 assign n_661 = ~(n_640 & in1_70_17_);
 assign n_660 = (in1_70_24_ | n_644);
 assign n_659 = ~(n_640 & in1_70_16_);
 assign n_658 = (in1_70_24_ | n_643);
 assign n_657 = ~(n_640 & in1_70_20_);
 assign n_656 = ~(in1_70_22_ & ~in1_70_24_);
 assign n_655 = ~(in1_68_22_ & in1_70_24_);
 assign n_654 = ~(in1_68_18_ & in1_70_24_);
 assign n_653 = ~(in1_70_19_ & ~in1_70_24_);
 assign n_652 = ~(n_640 & in1_70_2_);
 assign n_651 = ~(n_640 & in1_70_14_);
 assign n_650 = ~(n_640 & in1_70_13_);
 assign n_649 = ~(in1_70_24_ & n_1599);
 assign n_648 = ~(in1_70_21_ & ~in1_70_24_);
 assign n_647 = (in1_70_24_ | n_639);
 assign n_646 = ~(n_640 & in1_70_0_);
 assign n_645 = ~(n_640 & in1_70_18_);
 assign n_644 = ~in1_70_10_;
 assign n_643 = ~in1_70_8_;
 assign n_642 = ~in1_70_1_;
 assign n_641 = ~in1_70_11_;
 assign n_640 = ~in1_70_24_;
 assign n_639 = ~in1_70_12_;
 assign n_638 = ~in1_70_5_;
 assign n_637 = ~in1_70_3_;
 assign n_636 = ~(in1_70_24_ & in1_68_1_);
 assign n_635 = ~(in1_70_24_ & in1_68_19_);
 assign n_634 = ~(in1_70_24_ & in1_68_15_);
 assign n_633 = ~(in1_70_24_ & in1_68_6_);
 assign n_632 = ~(in1_70_7_ & ~in1_70_24_);
 assign n_631 = ~(in1_70_24_ & in1_68_20_);
 assign n_630 = ~(in1_70_6_ & ~in1_70_24_);
 assign n_629 = ~(in1_70_24_ & in1_68_0_);
 assign n_628 = ~(in1_70_24_ & in1_68_13_);
 assign n_627 = ~(in1_70_4_ & ~in1_70_24_);
 assign n_626 = ~(in1_70_24_ & in1_68_2_);
 assign n_625 = ~(in1_70_9_ & ~in1_70_24_);
 assign n_624 = ~(in1_70_24_ & in1_68_7_);
 assign n_623 = ~(in1_70_24_ & in1_68_3_);
 assign n_622 = ~(in1_70_24_ & in1_68_11_);
 assign n_621 = ~(in1_70_24_ & in1_68_10_);
 assign n_620 = ~(in1_70_24_ & in1_68_9_);
 assign n_619 = ~(in1_70_24_ & in1_68_21_);
 assign n_618 = ~(in1_70_24_ & in1_68_5_);
 assign n_617 = ~(in1_70_24_ & in1_68_4_);
 assign n_616 = ~(in1_70_24_ & in1_68_8_);
 assign n_615 = ~(in1_70_24_ & in1_68_14_);
 assign n_614 = ~(in1_70_24_ & in1_68_12_);
 assign in1_2_0_ = ~(n_613 & (in1_1_24_ | n_612));
 assign n_613 = ~(in1_1_24_ & {in1[48]});
 assign n_612 = ~in1_1_0_;
 assign in1_74_8_ = ~(n_604 & n_605);
 assign in1_74_20_ = ~(n_603 & n_581);
 assign in1_74_17_ = ~(n_609 & n_610);
 assign in1_74_10_ = ~(n_608 & n_565);
 assign in1_74_16_ = ~(n_580 & ~(n_587 & in1_73_16_));
 assign in1_74_9_ = ~(n_607 & n_561);
 assign in1_74_23_ = ~(n_597 & n_606);
 assign in1_74_19_ = ~(n_572 & ~(n_587 & in1_73_19_));
 assign in1_74_15_ = ~(n_602 & n_560);
 assign in1_74_7_ = ~(n_576 & n_578);
 assign in1_74_6_ = ~(n_574 & n_563);
 assign in1_74_14_ = ~(n_599 & n_571);
 assign in1_74_13_ = ~(n_596 & n_559);
 assign in1_74_22_ = ~(n_564 & ~(n_587 & in1_73_22_));
 assign in1_74_21_ = ~(n_575 & ~(n_587 & in1_73_21_));
 assign in1_74_4_ = ~(n_600 & n_568);
 assign in1_74_3_ = ~(n_598 & n_570);
 assign in1_74_18_ = ~(n_592 & n_579);
 assign in1_74_5_ = ~(n_569 & n_562);
 assign in1_74_2_ = ~(n_601 & n_582);
 assign in1_74_12_ = ~(n_594 & n_567);
 assign in1_74_1_ = ~(n_577 & n_573);
 assign in1_74_0_ = ~(n_593 & n_595);
 assign in1_74_11_ = ~(n_611 & n_566);
 assign n_611 = (in1_73_24_ | n_590);
 assign n_610 = ~(in1_71_16_ & in1_73_24_);
 assign n_609 = ~(n_587 & in1_73_17_);
 assign n_608 = (in1_73_24_ | n_591);
 assign n_607 = ~(n_587 & in1_73_9_);
 assign n_606 = ~(in1_71_22_ & in1_73_24_);
 assign n_605 = ~(in1_71_7_ & in1_73_24_);
 assign n_604 = ~(n_587 & in1_73_8_);
 assign n_603 = (in1_73_24_ | n_584);
 assign n_602 = (in1_73_24_ | n_583);
 assign n_601 = ~(n_587 & in1_73_2_);
 assign n_600 = (in1_73_24_ | n_589);
 assign n_599 = (in1_73_24_ | n_588);
 assign n_598 = ~(n_587 & in1_73_3_);
 assign n_597 = ~(in1_73_23_ & ~in1_73_24_);
 assign n_596 = (in1_73_24_ | n_585);
 assign n_595 = ~(in1_73_24_ & n_1572);
 assign n_594 = (in1_73_24_ | n_586);
 assign n_593 = ~(n_587 & in1_73_0_);
 assign n_592 = ~(n_587 & in1_73_18_);
 assign n_591 = ~in1_73_10_;
 assign n_590 = ~in1_73_11_;
 assign n_589 = ~in1_73_4_;
 assign n_588 = ~in1_73_14_;
 assign n_587 = ~in1_73_24_;
 assign n_586 = ~in1_73_12_;
 assign n_585 = ~in1_73_13_;
 assign n_584 = ~in1_73_20_;
 assign n_583 = ~in1_73_15_;
 assign n_582 = ~(in1_73_24_ & in1_71_1_);
 assign n_581 = ~(in1_73_24_ & in1_71_19_);
 assign n_580 = ~(in1_73_24_ & in1_71_15_);
 assign n_579 = ~(in1_73_24_ & in1_71_17_);
 assign n_578 = ~(in1_73_24_ & in1_71_6_);
 assign n_577 = ~(in1_73_1_ & ~in1_73_24_);
 assign n_576 = ~(in1_73_7_ & ~in1_73_24_);
 assign n_575 = ~(in1_73_24_ & in1_71_20_);
 assign n_574 = ~(in1_73_6_ & ~in1_73_24_);
 assign n_573 = ~(in1_73_24_ & in1_71_0_);
 assign n_572 = ~(in1_73_24_ & in1_71_18_);
 assign n_571 = ~(in1_73_24_ & in1_71_13_);
 assign n_570 = ~(in1_73_24_ & in1_71_2_);
 assign n_569 = ~(in1_73_5_ & ~in1_73_24_);
 assign n_568 = ~(in1_73_24_ & in1_71_3_);
 assign n_567 = ~(in1_73_24_ & in1_71_11_);
 assign n_566 = ~(in1_73_24_ & in1_71_10_);
 assign n_565 = ~(in1_73_24_ & in1_71_9_);
 assign n_564 = ~(in1_73_24_ & in1_71_21_);
 assign n_563 = ~(in1_73_24_ & in1_71_5_);
 assign n_562 = ~(in1_73_24_ & in1_71_4_);
 assign n_561 = ~(in1_73_24_ & in1_71_8_);
 assign n_560 = ~(in1_73_24_ & in1_71_14_);
 assign n_559 = ~(in1_73_24_ & in1_71_12_);
 assign in1_77_8_ = ~(n_547 & n_549);
 assign in1_77_20_ = ~(n_525 & ~(n_528 & in1_76_20_));
 assign in1_77_17_ = ~(n_554 & n_556);
 assign in1_77_10_ = ~(n_552 & n_553);
 assign in1_77_16_ = ~(n_548 & n_524);
 assign in1_77_9_ = ~(n_551 & n_514);
 assign in1_77_23_ = ~(n_529 & n_550);
 assign in1_77_19_ = ~(n_540 & n_541);
 assign in1_77_15_ = ~(n_544 & n_558);
 assign in1_77_7_ = ~(n_546 & n_522);
 assign in1_77_6_ = ~(n_543 & n_516);
 assign in1_77_14_ = ~(n_537 & n_520);
 assign in1_77_13_ = ~(n_513 & ~(n_528 & in1_76_13_));
 assign in1_77_22_ = ~(n_545 & n_557);
 assign in1_77_21_ = ~(n_533 & n_535);
 assign in1_77_4_ = ~(n_538 & n_518);
 assign in1_77_3_ = ~(n_536 & n_519);
 assign in1_77_18_ = ~(n_542 & n_523);
 assign in1_77_5_ = ~(n_555 & n_515);
 assign in1_77_2_ = ~(n_539 & n_526);
 assign in1_77_12_ = ~(n_530 & n_531);
 assign in1_77_1_ = ~(n_532 & n_521);
 assign in1_77_0_ = ~(n_512 & n_534);
 assign in1_77_11_ = ~(n_517 & ~(n_528 & in1_76_11_));
 assign n_558 = ~(in1_74_14_ & in1_76_24_);
 assign n_557 = ~(in1_74_21_ & in1_76_24_);
 assign n_556 = ~(in1_74_16_ & in1_76_24_);
 assign n_555 = ~(n_528 & in1_76_5_);
 assign n_554 = ~(n_528 & in1_76_17_);
 assign n_553 = ~(in1_74_9_ & in1_76_24_);
 assign n_552 = ~(n_528 & in1_76_10_);
 assign n_551 = (in1_76_24_ | n_527);
 assign n_550 = ~(in1_74_22_ & in1_76_24_);
 assign n_549 = ~(in1_74_7_ & in1_76_24_);
 assign n_548 = ~(n_528 & in1_76_16_);
 assign n_547 = ~(n_528 & in1_76_8_);
 assign n_546 = ~(n_528 & in1_76_7_);
 assign n_545 = ~(in1_76_22_ & ~in1_76_24_);
 assign n_544 = ~(in1_76_15_ & ~in1_76_24_);
 assign n_543 = ~(n_528 & in1_76_6_);
 assign n_542 = ~(n_528 & in1_76_18_);
 assign n_541 = ~(in1_74_18_ & in1_76_24_);
 assign n_540 = ~(in1_76_19_ & ~in1_76_24_);
 assign n_539 = ~(n_528 & in1_76_2_);
 assign n_538 = ~(n_528 & in1_76_4_);
 assign n_537 = ~(n_528 & in1_76_14_);
 assign n_536 = ~(n_528 & in1_76_3_);
 assign n_535 = ~(in1_74_20_ & in1_76_24_);
 assign n_534 = ~(in1_76_24_ & n_1542);
 assign n_533 = ~(in1_76_21_ & ~in1_76_24_);
 assign n_532 = ~(n_528 & in1_76_1_);
 assign n_531 = ~(in1_74_11_ & in1_76_24_);
 assign n_530 = ~(n_528 & in1_76_12_);
 assign n_529 = ~(in1_76_23_ & ~in1_76_24_);
 assign n_528 = ~in1_76_24_;
 assign n_527 = ~in1_76_9_;
 assign n_526 = ~(in1_76_24_ & in1_74_1_);
 assign n_525 = ~(in1_76_24_ & in1_74_19_);
 assign n_524 = ~(in1_76_24_ & in1_74_15_);
 assign n_523 = ~(in1_76_24_ & in1_74_17_);
 assign n_522 = ~(in1_76_24_ & in1_74_6_);
 assign n_521 = ~(in1_76_24_ & in1_74_0_);
 assign n_520 = ~(in1_76_24_ & in1_74_13_);
 assign n_519 = ~(in1_76_24_ & in1_74_2_);
 assign n_518 = ~(in1_76_24_ & in1_74_3_);
 assign n_517 = ~(in1_76_24_ & in1_74_10_);
 assign n_516 = ~(in1_76_24_ & in1_74_5_);
 assign n_515 = ~(in1_76_24_ & in1_74_4_);
 assign n_514 = ~(in1_76_24_ & in1_74_8_);
 assign n_513 = ~(in1_76_24_ & in1_74_12_);
 assign n_512 = ~(in1_76_0_ & ~in1_76_24_);
 assign in1_80_8_ = ~(n_501 & ~(n_471 & in1_79_8_));
 assign in1_80_20_ = ~(n_499 & n_505);
 assign in1_80_17_ = ~(n_507 & n_508);
 assign in1_80_10_ = ~(n_506 & n_465);
 assign in1_80_16_ = ~(n_500 & n_503);
 assign in1_80_9_ = ~(n_504 & n_464);
 assign in1_80_23_ = ~(n_511 & n_494);
 assign in1_80_19_ = ~(n_493 & ~(n_471 & in1_79_19_));
 assign in1_80_15_ = ~(n_502 & ~(n_471 & in1_79_15_));
 assign in1_80_7_ = ~(n_497 & n_498);
 assign in1_80_6_ = ~(n_495 & ~(n_471 & in1_79_6_));
 assign in1_80_14_ = ~(n_488 & n_492);
 assign in1_80_13_ = ~(n_482 & n_486);
 assign in1_80_22_ = ~(n_496 & n_509);
 assign in1_80_21_ = ~(n_479 & n_485);
 assign in1_80_4_ = ~(n_489 & n_491);
 assign in1_80_3_ = ~(n_487 & n_481);
 assign in1_80_18_ = ~(n_473 & n_478);
 assign in1_80_5_ = ~(n_483 & ~(n_471 & in1_79_5_));
 assign in1_80_2_ = ~(n_490 & n_467);
 assign in1_80_12_ = ~(n_475 & n_476);
 assign in1_80_1_ = ~(n_477 & n_466);
 assign in1_80_0_ = ~(n_474 & n_480);
 assign in1_80_11_ = ~(n_510 & n_484);
 assign n_511 = ~(in1_79_23_ & ~in1_79_24_);
 assign n_510 = ~(n_471 & in1_79_11_);
 assign n_509 = ~(in1_77_21_ & in1_79_24_);
 assign n_508 = ~(in1_77_16_ & in1_79_24_);
 assign n_507 = ~(n_471 & in1_79_17_);
 assign n_506 = ~(n_471 & in1_79_10_);
 assign n_505 = ~(in1_77_19_ & in1_79_24_);
 assign n_504 = ~(n_471 & in1_79_9_);
 assign n_503 = ~(in1_77_15_ & in1_79_24_);
 assign n_502 = ~(in1_77_14_ & in1_79_24_);
 assign n_501 = ~(in1_77_7_ & in1_79_24_);
 assign n_500 = (in1_79_24_ | n_469);
 assign n_499 = ~(in1_79_20_ & ~in1_79_24_);
 assign n_498 = ~(in1_77_6_ & in1_79_24_);
 assign n_497 = ~(n_471 & in1_79_7_);
 assign n_496 = ~(in1_79_22_ & ~in1_79_24_);
 assign n_495 = ~(in1_77_5_ & in1_79_24_);
 assign n_494 = ~(in1_77_22_ & in1_79_24_);
 assign n_493 = ~(in1_77_18_ & in1_79_24_);
 assign n_492 = ~(in1_77_13_ & in1_79_24_);
 assign n_491 = ~(in1_77_3_ & in1_79_24_);
 assign n_490 = ~(n_471 & in1_79_2_);
 assign n_489 = ~(n_471 & in1_79_4_);
 assign n_488 = (in1_79_24_ | n_472);
 assign n_487 = ~(n_471 & in1_79_3_);
 assign n_486 = ~(in1_77_12_ & in1_79_24_);
 assign n_485 = ~(in1_77_20_ & in1_79_24_);
 assign n_484 = ~(in1_77_10_ & in1_79_24_);
 assign n_483 = ~(in1_77_4_ & in1_79_24_);
 assign n_482 = ~(n_471 & in1_79_13_);
 assign n_481 = ~(in1_77_2_ & in1_79_24_);
 assign n_480 = ~(in1_79_24_ & n_1585);
 assign n_479 = ~(in1_79_21_ & ~in1_79_24_);
 assign n_478 = ~(in1_77_17_ & in1_79_24_);
 assign n_477 = ~(n_471 & in1_79_1_);
 assign n_476 = ~(in1_77_11_ & in1_79_24_);
 assign n_475 = (in1_79_24_ | n_470);
 assign n_474 = (in1_79_24_ | n_468);
 assign n_473 = ~(n_471 & in1_79_18_);
 assign n_472 = ~in1_79_14_;
 assign n_471 = ~in1_79_24_;
 assign n_470 = ~in1_79_12_;
 assign n_469 = ~in1_79_16_;
 assign n_468 = ~in1_79_0_;
 assign n_467 = ~(in1_79_24_ & in1_77_1_);
 assign n_466 = ~(in1_79_24_ & in1_77_0_);
 assign n_465 = ~(in1_79_24_ & in1_77_9_);
 assign n_464 = ~(in1_79_24_ & in1_77_8_);
 assign in1_83_8_ = ~(n_456 & ~(n_434 & in1_82_8_));
 assign in1_83_20_ = ~(n_455 & ~(in1_80_19_ & in1_82_24_));
 assign in1_83_17_ = ~(n_461 & ~(n_434 & in1_82_17_));
 assign in1_83_10_ = ~(n_460 & ~(in1_80_9_ & in1_82_24_));
 assign in1_83_16_ = ~(n_458 & ~(n_434 & in1_82_16_));
 assign in1_83_9_ = ~(n_459 & ~(in1_80_8_ & in1_82_24_));
 assign in1_83_23_ = ~(n_450 & ~(n_434 & in1_82_23_));
 assign in1_83_19_ = ~(n_442 & ~(in1_80_18_ & in1_82_24_));
 assign in1_83_15_ = ~(n_452 & n_457);
 assign in1_83_7_ = ~(n_454 & ~(in1_80_6_ & in1_82_24_));
 assign in1_83_6_ = ~(n_451 & ~(n_434 & in1_82_6_));
 assign in1_83_14_ = ~(n_448 & ~(n_434 & in1_82_14_));
 assign in1_83_13_ = ~(n_444 & ~(n_434 & in1_82_13_));
 assign in1_83_22_ = ~(n_453 & n_462);
 assign in1_83_21_ = ~(n_439 & n_443);
 assign in1_83_4_ = ~(n_447 & ~(n_434 & in1_82_4_));
 assign in1_83_3_ = ~(n_445 & ~(in1_80_2_ & in1_82_24_));
 assign in1_83_18_ = ~(n_438 & ~(n_434 & in1_82_18_));
 assign in1_83_5_ = ~(n_463 & ~(n_434 & in1_82_5_));
 assign in1_83_2_ = ~(n_446 & n_441);
 assign in1_83_12_ = ~(n_436 & ~(n_434 & in1_82_12_));
 assign in1_83_1_ = ~(n_437 & ~(in1_80_0_ & in1_82_24_));
 assign in1_83_0_ = ~(n_435 & n_440);
 assign in1_83_11_ = ~(n_449 & ~(n_434 & in1_82_11_));
 assign n_463 = ~(in1_80_4_ & in1_82_24_);
 assign n_462 = ~(in1_80_21_ & in1_82_24_);
 assign n_461 = ~(in1_80_16_ & in1_82_24_);
 assign n_460 = ~(n_434 & in1_82_10_);
 assign n_459 = ~(n_434 & in1_82_9_);
 assign n_458 = ~(in1_80_15_ & in1_82_24_);
 assign n_457 = ~(in1_80_14_ & in1_82_24_);
 assign n_456 = ~(in1_80_7_ & in1_82_24_);
 assign n_455 = ~(n_434 & in1_82_20_);
 assign n_454 = ~(n_434 & in1_82_7_);
 assign n_453 = ~(in1_82_22_ & ~in1_82_24_);
 assign n_452 = ~(in1_82_15_ & ~in1_82_24_);
 assign n_451 = ~(in1_80_5_ & in1_82_24_);
 assign n_450 = ~(in1_80_22_ & in1_82_24_);
 assign n_449 = ~(in1_80_10_ & in1_82_24_);
 assign n_448 = ~(in1_80_13_ & in1_82_24_);
 assign n_447 = ~(in1_80_3_ & in1_82_24_);
 assign n_446 = ~(n_434 & in1_82_2_);
 assign n_445 = ~(n_434 & in1_82_3_);
 assign n_444 = ~(in1_80_12_ & in1_82_24_);
 assign n_443 = ~(in1_80_20_ & in1_82_24_);
 assign n_442 = ~(in1_82_19_ & ~in1_82_24_);
 assign n_441 = ~(in1_80_1_ & in1_82_24_);
 assign n_440 = ~(in1_82_24_ & n_1588);
 assign n_439 = ~(in1_82_21_ & ~in1_82_24_);
 assign n_438 = ~(in1_80_17_ & in1_82_24_);
 assign n_437 = ~(n_434 & in1_82_1_);
 assign n_436 = ~(in1_80_11_ & in1_82_24_);
 assign n_435 = ~(n_434 & in1_82_0_);
 assign n_434 = ~in1_82_24_;
 assign in1_86_8_ = ~(n_424 & ~(n_407 & in1_85_8_));
 assign in1_86_20_ = ~(n_428 & ~(n_407 & in1_85_20_));
 assign in1_86_17_ = ~(n_430 & ~(n_407 & in1_85_17_));
 assign in1_86_10_ = ~(n_429 & ~(n_407 & in1_85_10_));
 assign in1_86_16_ = ~(n_426 & ~(n_407 & in1_85_16_));
 assign in1_86_9_ = ~(n_433 & ~(in1_83_8_ & in1_85_24_));
 assign in1_86_23_ = ~(n_427 & ~(n_407 & in1_85_23_));
 assign in1_86_19_ = ~(n_419 & ~(n_407 & in1_85_19_));
 assign in1_86_15_ = ~(n_422 & n_425);
 assign in1_86_7_ = ~(n_423 & (in1_85_24_ | n_408));
 assign in1_86_6_ = ~(n_421 & ~(n_407 & in1_85_6_));
 assign in1_86_14_ = ~(n_417 & n_418);
 assign in1_86_13_ = ~(n_415 & (in1_85_24_ | n_406));
 assign in1_86_22_ = ~(n_431 & ~(n_407 & in1_85_22_));
 assign in1_86_21_ = ~(n_414 & ~(n_407 & in1_85_21_));
 assign in1_86_4_ = ((in1_85_4_ & ~in1_85_24_) | (in1_83_3_ & in1_85_24_));
 assign in1_86_3_ = ~(n_416 & ~(in1_83_2_ & in1_85_24_));
 assign in1_86_18_ = ~(n_412 & ~(n_407 & in1_85_18_));
 assign in1_86_5_ = ~(n_420 & ~(n_407 & in1_85_5_));
 assign in1_86_2_ = ((in1_85_2_ & ~in1_85_24_) | (in1_83_1_ & in1_85_24_));
 assign in1_86_12_ = ~(n_410 & ~(n_407 & in1_85_12_));
 assign in1_86_1_ = ~(n_411 & ~(in1_83_0_ & in1_85_24_));
 assign in1_86_0_ = ~(n_409 & n_413);
 assign in1_86_11_ = ~(n_432 & ~(in1_83_10_ & in1_85_24_));
 assign n_433 = ~(n_407 & in1_85_9_);
 assign n_432 = ~(n_407 & in1_85_11_);
 assign n_431 = ~(in1_83_21_ & in1_85_24_);
 assign n_430 = ~(in1_83_16_ & in1_85_24_);
 assign n_429 = ~(in1_83_9_ & in1_85_24_);
 assign n_428 = ~(in1_83_19_ & in1_85_24_);
 assign n_427 = ~(in1_83_22_ & in1_85_24_);
 assign n_426 = ~(in1_83_15_ & in1_85_24_);
 assign n_425 = ~(in1_83_14_ & in1_85_24_);
 assign n_424 = ~(in1_83_7_ & in1_85_24_);
 assign n_423 = ~(in1_83_6_ & in1_85_24_);
 assign n_422 = ~(n_407 & in1_85_15_);
 assign n_421 = ~(in1_83_5_ & in1_85_24_);
 assign n_420 = ~(in1_83_4_ & in1_85_24_);
 assign n_419 = ~(in1_83_18_ & in1_85_24_);
 assign n_418 = ~(in1_83_13_ & in1_85_24_);
 assign n_417 = ~(n_407 & in1_85_14_);
 assign n_416 = ~(n_407 & in1_85_3_);
 assign n_415 = ~(in1_83_12_ & in1_85_24_);
 assign n_414 = ~(in1_83_20_ & in1_85_24_);
 assign n_413 = ~(in1_85_24_ & n_1561);
 assign n_412 = ~(in1_83_17_ & in1_85_24_);
 assign n_411 = ~(n_407 & in1_85_1_);
 assign n_410 = ~(in1_83_11_ & in1_85_24_);
 assign n_409 = ~(n_407 & in1_85_0_);
 assign n_408 = ~in1_85_7_;
 assign n_407 = ~in1_85_24_;
 assign n_406 = ~in1_85_13_;
 assign in1_89_8_ = ~(n_396 & ~(n_377 & in1_88_8_));
 assign in1_89_20_ = ~(n_400 & ~(n_377 & in1_88_20_));
 assign in1_89_17_ = ~(n_403 & ~(n_377 & in1_88_17_));
 assign in1_89_10_ = ~(n_401 & ~(n_377 & in1_88_10_));
 assign in1_89_16_ = ~(n_398 & ~(n_377 & in1_88_16_));
 assign in1_89_9_ = ~(n_399 & ~(n_377 & in1_88_9_));
 assign in1_89_23_ = ~(n_405 & n_392);
 assign in1_89_19_ = ~(n_389 & n_390);
 assign in1_89_15_ = ~(n_397 & ~(n_377 & in1_88_15_));
 assign in1_89_7_ = ~(n_395 & ~(n_377 & in1_88_7_));
 assign in1_89_6_ = ~(n_393 & ~(n_377 & in1_88_6_));
 assign in1_89_14_ = ~(n_388 & ~(n_377 & in1_88_14_));
 assign in1_89_13_ = ~(n_385 & ~(n_377 & in1_88_13_));
 assign in1_89_22_ = ~(n_394 & n_404);
 assign in1_89_21_ = ~(n_384 & ~(n_377 & in1_88_21_));
 assign in1_89_4_ = ~(n_387 & ~(n_377 & in1_88_4_));
 assign in1_89_3_ = ~(n_386 & ~(in1_86_2_ & in1_88_24_));
 assign in1_89_18_ = ~(n_381 & ~(n_377 & in1_88_18_));
 assign in1_89_5_ = ~(n_402 & n_378);
 assign in1_89_2_ = ~(n_382 & ~(n_377 & in1_88_2_));
 assign in1_89_12_ = ~(n_379 & ~(n_377 & in1_88_12_));
 assign in1_89_1_ = ~(n_380 & ~(in1_86_0_ & in1_88_24_));
 assign in1_89_0_ = ~(n_391 & ~(in1_88_24_ & n_1584));
 assign in1_89_11_ = ~(n_383 & ~(n_377 & in1_88_11_));
 assign n_405 = ~(in1_88_23_ & ~in1_88_24_);
 assign n_404 = ~(in1_86_21_ & in1_88_24_);
 assign n_403 = ~(in1_86_16_ & in1_88_24_);
 assign n_402 = ~(n_377 & in1_88_5_);
 assign n_401 = ~(in1_86_9_ & in1_88_24_);
 assign n_400 = ~(in1_86_19_ & in1_88_24_);
 assign n_399 = ~(in1_86_8_ & in1_88_24_);
 assign n_398 = ~(in1_86_15_ & in1_88_24_);
 assign n_397 = ~(in1_86_14_ & in1_88_24_);
 assign n_396 = ~(in1_86_7_ & in1_88_24_);
 assign n_395 = ~(in1_86_6_ & in1_88_24_);
 assign n_394 = ~(in1_88_22_ & ~in1_88_24_);
 assign n_393 = ~(in1_86_5_ & in1_88_24_);
 assign n_392 = ~(in1_86_22_ & in1_88_24_);
 assign n_391 = ~(n_377 & in1_88_0_);
 assign n_390 = ~(in1_86_18_ & in1_88_24_);
 assign n_389 = ~(in1_88_19_ & ~in1_88_24_);
 assign n_388 = ~(in1_86_13_ & in1_88_24_);
 assign n_387 = ~(in1_86_3_ & in1_88_24_);
 assign n_386 = ~(n_377 & in1_88_3_);
 assign n_385 = ~(in1_86_12_ & in1_88_24_);
 assign n_384 = ~(in1_86_20_ & in1_88_24_);
 assign n_383 = ~(in1_86_10_ & in1_88_24_);
 assign n_382 = ~(in1_86_1_ & in1_88_24_);
 assign n_381 = ~(in1_86_17_ & in1_88_24_);
 assign n_380 = ~(n_377 & in1_88_1_);
 assign n_379 = ~(in1_86_11_ & in1_88_24_);
 assign n_378 = ~(in1_86_4_ & in1_88_24_);
 assign n_377 = ~in1_88_24_;
 assign asc001_0_8_ = ~in1_121_24_;
 assign asc001_0_1_ = ~in1_142_24_;
 assign asc001_0_2_ = ~in1_139_24_;
 assign asc001_0_3_ = ~in1_136_24_;
 assign asc001_0_4_ = ~in1_133_24_;
 assign asc001_0_5_ = ~in1_130_24_;
 assign asc001_0_6_ = ~in1_127_24_;
 assign asc001_0_7_ = ~in1_124_24_;
 assign asc001_0_36_ = ~in1_37_24_;
 assign asc001_0_9_ = ~in1_118_24_;
 assign asc001_0_10_ = ~in1_115_24_;
 assign asc001_0_11_ = ~in1_112_24_;
 assign asc001_0_12_ = ~in1_109_24_;
 assign asc001_0_13_ = ~n_1440;
 assign asc001_0_14_ = ~n_1438;
 assign asc001_0_15_ = ~n_1407;
 assign asc001_0_16_ = ~n_1413;
 assign asc001_0_26_ = ~in1_67_24_;
 assign asc001_0_18_ = ~n_1415;
 assign asc001_0_19_ = ~n_1408;
 assign asc001_0_20_ = ~n_1406;
 assign asc001_0_21_ = ~n_1462;
 assign asc001_0_22_ = ~in1_79_24_;
 assign asc001_0_23_ = ~n_1461;
 assign asc001_0_24_ = ~in1_73_24_;
 assign asc001_0_25_ = ~in1_70_24_;
 assign asc001_0_17_ = ~n_1414;
 assign asc001_0_27_ = ~in1_64_24_;
 assign asc001_0_28_ = ~n_1494;
 assign asc001_0_29_ = ~n_1492;
 assign asc001_0_30_ = ~in1_55_24_;
 assign asc001_0_31_ = ~in1_52_24_;
 assign asc001_0_32_ = ~n_1487;
 assign asc001_0_33_ = ~in1_46_24_;
 assign asc001_0_34_ = ~n_1485;
 assign asc001_0_35_ = ~in1_40_24_;
 assign in1_92_8_ = ~(n_367 & ~(n_349 & in1_91_8_));
 assign in1_92_20_ = ~(n_371 & ~(n_349 & in1_91_20_));
 assign in1_92_17_ = ~(n_374 & ~(n_349 & in1_91_17_));
 assign in1_92_10_ = ~(n_372 & n_373);
 assign in1_92_16_ = ~(n_366 & ~(in1_89_15_ & in1_91_24_));
 assign in1_92_9_ = ~(n_369 & n_370);
 assign in1_92_23_ = ~(n_376 & ~(n_349 & in1_91_23_));
 assign in1_92_19_ = ~(n_361 & ~(n_349 & in1_91_19_));
 assign in1_92_15_ = ~(n_368 & ~(n_349 & in1_91_15_));
 assign in1_92_7_ = ~(n_365 & ~(in1_89_6_ & in1_91_24_));
 assign in1_92_6_ = ~(n_350 & ~(n_349 & in1_91_6_));
 assign in1_92_14_ = ~(n_360 & ~(n_349 & in1_91_14_));
 assign in1_92_13_ = ~(n_357 & ~(n_349 & in1_91_13_));
 assign in1_92_22_ = ~(n_375 & ~(n_349 & in1_91_22_));
 assign in1_92_21_ = ~(n_356 & ~(n_349 & in1_91_21_));
 assign in1_92_4_ = ~(n_359 & ~(n_349 & in1_91_4_));
 assign in1_92_3_ = ~(n_358 & ~(in1_89_2_ & in1_91_24_));
 assign in1_92_18_ = ~(n_353 & ~(n_349 & in1_91_18_));
 assign in1_92_5_ = ~(n_362 & ~(n_349 & in1_91_5_));
 assign in1_92_2_ = ~(n_354 & ~(n_349 & in1_91_2_));
 assign in1_92_12_ = ~(n_351 & ~(in1_89_11_ & in1_91_24_));
 assign in1_92_1_ = ~(n_352 & n_364);
 assign in1_92_0_ = ~(n_363 & ~(in1_91_24_ & n_1532));
 assign in1_92_11_ = ~(n_355 & ~(n_349 & in1_91_11_));
 assign n_376 = ~(in1_89_22_ & in1_91_24_);
 assign n_375 = ~(in1_89_21_ & in1_91_24_);
 assign n_374 = ~(in1_89_16_ & in1_91_24_);
 assign n_373 = ~(in1_89_9_ & in1_91_24_);
 assign n_372 = ~(n_349 & in1_91_10_);
 assign n_371 = ~(in1_89_19_ & in1_91_24_);
 assign n_370 = ~(in1_89_8_ & in1_91_24_);
 assign n_369 = ~(n_349 & in1_91_9_);
 assign n_368 = ~(in1_89_14_ & in1_91_24_);
 assign n_367 = ~(in1_89_7_ & in1_91_24_);
 assign n_366 = ~(n_349 & in1_91_16_);
 assign n_365 = ~(n_349 & in1_91_7_);
 assign n_364 = ~(in1_89_0_ & in1_91_24_);
 assign n_363 = ~(n_349 & in1_91_0_);
 assign n_362 = ~(in1_89_4_ & in1_91_24_);
 assign n_361 = ~(in1_89_18_ & in1_91_24_);
 assign n_360 = ~(in1_89_13_ & in1_91_24_);
 assign n_359 = ~(in1_89_3_ & in1_91_24_);
 assign n_358 = ~(n_349 & in1_91_3_);
 assign n_357 = ~(in1_89_12_ & in1_91_24_);
 assign n_356 = ~(in1_89_20_ & in1_91_24_);
 assign n_355 = ~(in1_89_10_ & in1_91_24_);
 assign n_354 = ~(in1_89_1_ & in1_91_24_);
 assign n_353 = ~(in1_89_17_ & in1_91_24_);
 assign n_352 = ~(n_349 & in1_91_1_);
 assign n_351 = ~(n_349 & in1_91_12_);
 assign n_350 = ~(in1_89_5_ & in1_91_24_);
 assign n_349 = ~in1_91_24_;
 assign in1_95_8_ = ~(n_339 & ~(n_316 & in1_94_8_));
 assign in1_95_20_ = ~(n_344 & ~(n_316 & in1_94_20_));
 assign in1_95_17_ = ~(n_346 & ~(n_316 & in1_94_17_));
 assign in1_95_10_ = ~(n_345 & ~(n_316 & in1_94_10_));
 assign in1_95_16_ = ~(n_341 & ~(n_316 & in1_94_16_));
 assign in1_95_9_ = ~(n_342 & n_343);
 assign in1_95_23_ = ~(n_333 & ~(n_316 & in1_94_23_));
 assign in1_95_19_ = ~(n_331 & n_317);
 assign in1_95_15_ = ~(n_340 & ~(n_316 & in1_94_15_));
 assign in1_95_7_ = ~(n_337 & n_338);
 assign in1_95_6_ = ~(n_334 & ~(n_316 & in1_94_6_));
 assign in1_95_14_ = ~(n_330 & ~(n_316 & in1_94_14_));
 assign in1_95_13_ = ~(n_327 & ~(n_316 & in1_94_13_));
 assign in1_95_22_ = ~(n_336 & n_347);
 assign in1_95_21_ = ~(n_321 & n_326);
 assign in1_95_4_ = ~(n_329 & ~(n_316 & in1_94_4_));
 assign in1_95_3_ = ~(n_323 & ~(n_316 & in1_94_3_));
 assign in1_95_18_ = ~(n_320 & ~(n_316 & in1_94_18_));
 assign in1_95_5_ = ~(n_348 & ~(n_316 & in1_94_5_));
 assign in1_95_2_ = ~(n_328 & n_324);
 assign in1_95_12_ = ~(n_318 & ~(n_316 & in1_94_12_));
 assign in1_95_1_ = ~(n_319 & n_335);
 assign in1_95_0_ = ~(n_332 & n_322);
 assign in1_95_11_ = ~(n_325 & ~(n_316 & in1_94_11_));
 assign n_348 = ~(in1_92_4_ & in1_94_24_);
 assign n_347 = ~(in1_92_21_ & in1_94_24_);
 assign n_346 = ~(in1_92_16_ & in1_94_24_);
 assign n_345 = ~(in1_92_9_ & in1_94_24_);
 assign n_344 = ~(in1_92_19_ & in1_94_24_);
 assign n_343 = ~(in1_92_8_ & in1_94_24_);
 assign n_342 = ~(n_316 & in1_94_9_);
 assign n_341 = ~(in1_92_15_ & in1_94_24_);
 assign n_340 = ~(in1_92_14_ & in1_94_24_);
 assign n_339 = ~(in1_92_7_ & in1_94_24_);
 assign n_338 = ~(in1_92_6_ & in1_94_24_);
 assign n_337 = ~(n_316 & in1_94_7_);
 assign n_336 = ~(in1_94_22_ & ~in1_94_24_);
 assign n_335 = ~(in1_92_0_ & in1_94_24_);
 assign n_334 = ~(in1_92_5_ & in1_94_24_);
 assign n_333 = ~(in1_92_22_ & in1_94_24_);
 assign n_332 = ~(n_316 & in1_94_0_);
 assign n_331 = ~(in1_94_19_ & ~in1_94_24_);
 assign n_330 = ~(in1_92_13_ & in1_94_24_);
 assign n_329 = ~(in1_92_3_ & in1_94_24_);
 assign n_328 = ~(n_316 & in1_94_2_);
 assign n_327 = ~(in1_92_12_ & in1_94_24_);
 assign n_326 = ~(in1_92_20_ & in1_94_24_);
 assign n_325 = ~(in1_92_10_ & in1_94_24_);
 assign n_324 = ~(in1_92_1_ & in1_94_24_);
 assign n_323 = ~(in1_92_2_ & in1_94_24_);
 assign n_322 = ~(in1_94_24_ & n_1557);
 assign n_321 = ~(in1_94_21_ & ~in1_94_24_);
 assign n_320 = ~(in1_92_17_ & in1_94_24_);
 assign n_319 = ~(n_316 & in1_94_1_);
 assign n_318 = ~(in1_92_11_ & in1_94_24_);
 assign n_317 = ~(in1_92_18_ & in1_94_24_);
 assign n_316 = ~in1_94_24_;
 assign in1_98_8_ = ~(n_307 & ~(n_290 & in1_97_8_));
 assign in1_98_20_ = ~(n_311 & ~(n_290 & in1_97_20_));
 assign in1_98_17_ = ~(n_313 & ~(in1_95_16_ & in1_97_24_));
 assign in1_98_10_ = ~(n_312 & ~(n_290 & in1_97_10_));
 assign in1_98_16_ = ~(n_315 & ~(n_290 & in1_97_16_));
 assign in1_98_9_ = ~(n_310 & ~(in1_95_8_ & in1_97_24_));
 assign in1_98_23_ = ~(n_309 & ~(n_290 & in1_97_23_));
 assign in1_98_19_ = ~(n_302 & ~(n_290 & in1_97_19_));
 assign in1_98_15_ = ~(n_305 & n_308);
 assign in1_98_7_ = ~(n_306 & ~(in1_95_6_ & in1_97_24_));
 assign in1_98_6_ = ~(n_304 & ~(n_290 & in1_97_6_));
 assign in1_98_14_ = ~(n_301 & ~(n_290 & in1_97_14_));
 assign in1_98_13_ = ~(n_298 & ~(n_290 & in1_97_13_));
 assign in1_98_22_ = ~(n_314 & ~(n_290 & in1_97_22_));
 assign in1_98_21_ = ~(n_297 & ~(n_290 & in1_97_21_));
 assign in1_98_4_ = ~(n_300 & ~(n_290 & in1_97_4_));
 assign in1_98_3_ = ~(n_299 & ~(in1_95_2_ & in1_97_24_));
 assign in1_98_18_ = ~(n_293 & ~(n_290 & in1_97_18_));
 assign in1_98_5_ = ~(n_303 & ~(n_290 & in1_97_5_));
 assign in1_98_2_ = ~(n_295 & ~(n_290 & in1_97_2_));
 assign in1_98_12_ = ~(n_291 & ~(n_290 & in1_97_12_));
 assign in1_98_1_ = ~(n_292 & ~(in1_95_0_ & in1_97_24_));
 assign in1_98_0_ = ~(n_294 & (in1_97_24_ | n_289));
 assign in1_98_11_ = ~(n_296 & ~(n_290 & in1_97_11_));
 assign n_315 = ~(in1_95_15_ & in1_97_24_);
 assign n_314 = ~(in1_95_21_ & in1_97_24_);
 assign n_313 = ~(n_290 & in1_97_17_);
 assign n_312 = ~(in1_95_9_ & in1_97_24_);
 assign n_311 = ~(in1_95_19_ & in1_97_24_);
 assign n_310 = ~(n_290 & in1_97_9_);
 assign n_309 = ~(in1_95_22_ & in1_97_24_);
 assign n_308 = ~(in1_95_14_ & in1_97_24_);
 assign n_307 = ~(in1_95_7_ & in1_97_24_);
 assign n_306 = ~(n_290 & in1_97_7_);
 assign n_305 = ~(in1_97_15_ & ~in1_97_24_);
 assign n_304 = ~(in1_95_5_ & in1_97_24_);
 assign n_303 = ~(in1_95_4_ & in1_97_24_);
 assign n_302 = ~(in1_95_18_ & in1_97_24_);
 assign n_301 = ~(in1_95_13_ & in1_97_24_);
 assign n_300 = ~(in1_95_3_ & in1_97_24_);
 assign n_299 = ~(n_290 & in1_97_3_);
 assign n_298 = ~(in1_95_12_ & in1_97_24_);
 assign n_297 = ~(in1_95_20_ & in1_97_24_);
 assign n_296 = ~(in1_95_10_ & in1_97_24_);
 assign n_295 = ~(in1_95_1_ & in1_97_24_);
 assign n_294 = ~(in1_97_24_ & n_1560);
 assign n_293 = ~(in1_95_17_ & in1_97_24_);
 assign n_292 = ~(n_290 & in1_97_1_);
 assign n_291 = ~(in1_95_11_ & in1_97_24_);
 assign n_290 = ~in1_97_24_;
 assign n_289 = ~in1_97_0_;
 assign in1_101_8_ = ~(n_279 & ~(n_261 & in1_100_8_));
 assign in1_101_20_ = ~(n_283 & ~(n_261 & in1_100_20_));
 assign in1_101_17_ = ~(n_286 & ~(n_261 & in1_100_17_));
 assign in1_101_10_ = ~(n_284 & ~(n_261 & in1_100_10_));
 assign in1_101_16_ = ~(n_278 & n_281);
 assign in1_101_9_ = ~(n_282 & ~(n_261 & in1_100_9_));
 assign in1_101_23_ = ~(n_288 & ~(n_261 & in1_100_23_));
 assign in1_101_19_ = ~(n_273 & ~(n_261 & in1_100_19_));
 assign in1_101_15_ = ~(n_262 & n_280);
 assign in1_101_7_ = ~(n_276 & n_277);
 assign in1_101_6_ = ~(n_274 & ~(n_261 & in1_100_6_));
 assign in1_101_14_ = ~(n_272 & ~(n_261 & in1_100_14_));
 assign in1_101_13_ = ~(n_269 & ~(n_261 & in1_100_13_));
 assign in1_101_22_ = ~(n_287 & ~(n_261 & in1_100_22_));
 assign in1_101_21_ = ~(n_268 & ~(n_261 & in1_100_21_));
 assign in1_101_4_ = ~(n_271 & ~(n_261 & in1_100_4_));
 assign in1_101_3_ = ~(n_266 & (in1_100_24_ | n_260));
 assign in1_101_18_ = ~(n_265 & ~(n_261 & in1_100_18_));
 assign in1_101_5_ = ~(n_285 & ~(in1_98_4_ & in1_100_24_));
 assign in1_101_2_ = ~(n_270 & ~(in1_98_1_ & in1_100_24_));
 assign in1_101_12_ = ~(n_263 & ~(n_261 & in1_100_12_));
 assign in1_101_1_ = ~(n_264 & ~(in1_98_0_ & in1_100_24_));
 assign in1_101_0_ = ~(n_275 & ~(in1_100_24_ & n_1564));
 assign in1_101_11_ = ~(n_267 & ~(n_261 & in1_100_11_));
 assign n_288 = ~(in1_98_22_ & in1_100_24_);
 assign n_287 = ~(in1_98_21_ & in1_100_24_);
 assign n_286 = ~(in1_98_16_ & in1_100_24_);
 assign n_285 = ~(n_261 & in1_100_5_);
 assign n_284 = ~(in1_98_9_ & in1_100_24_);
 assign n_283 = ~(in1_98_19_ & in1_100_24_);
 assign n_282 = ~(in1_98_8_ & in1_100_24_);
 assign n_281 = ~(in1_98_15_ & in1_100_24_);
 assign n_280 = ~(in1_98_14_ & in1_100_24_);
 assign n_279 = ~(in1_98_7_ & in1_100_24_);
 assign n_278 = ~(n_261 & in1_100_16_);
 assign n_277 = ~(in1_98_6_ & in1_100_24_);
 assign n_276 = ~(n_261 & in1_100_7_);
 assign n_275 = ~(n_261 & in1_100_0_);
 assign n_274 = ~(in1_98_5_ & in1_100_24_);
 assign n_273 = ~(in1_98_18_ & in1_100_24_);
 assign n_272 = ~(in1_98_13_ & in1_100_24_);
 assign n_271 = ~(in1_98_3_ & in1_100_24_);
 assign n_270 = ~(n_261 & in1_100_2_);
 assign n_269 = ~(in1_98_12_ & in1_100_24_);
 assign n_268 = ~(in1_98_20_ & in1_100_24_);
 assign n_267 = ~(in1_98_10_ & in1_100_24_);
 assign n_266 = ~(in1_98_2_ & in1_100_24_);
 assign n_265 = ~(in1_98_17_ & in1_100_24_);
 assign n_264 = ~(n_261 & in1_100_1_);
 assign n_263 = ~(in1_98_11_ & in1_100_24_);
 assign n_262 = ~(in1_100_15_ & ~in1_100_24_);
 assign n_261 = ~in1_100_24_;
 assign n_260 = ~in1_100_3_;
 assign in1_104_8_ = ~(n_249 & ~(n_230 & in1_103_8_));
 assign in1_104_20_ = ~(n_253 & ~(n_230 & in1_103_20_));
 assign in1_104_17_ = ~(n_256 & ~(n_230 & in1_103_17_));
 assign in1_104_10_ = ~(n_254 & n_255);
 assign in1_104_16_ = ~(n_251 & ~(n_230 & in1_103_16_));
 assign in1_104_9_ = ~(n_252 & ~(n_230 & in1_103_9_));
 assign in1_104_23_ = ~(n_246 & ~(n_230 & in1_103_23_));
 assign in1_104_19_ = ~(n_244 & ~(n_230 & in1_103_19_));
 assign in1_104_15_ = ~(n_250 & ~(n_230 & in1_103_15_));
 assign in1_104_7_ = ~(n_247 & n_248);
 assign in1_104_6_ = ~(n_259 & ~(n_230 & in1_103_6_));
 assign in1_104_14_ = ~(n_243 & ~(n_230 & in1_103_14_));
 assign in1_104_13_ = ~(n_239 & ~(n_230 & in1_103_13_));
 assign in1_104_22_ = ~(n_257 & ~(n_230 & in1_103_22_));
 assign in1_104_21_ = ~(n_234 & n_245);
 assign in1_104_4_ = ~(n_242 & ~(n_230 & in1_103_4_));
 assign in1_104_3_ = ~(n_240 & ~(in1_101_2_ & in1_103_24_));
 assign in1_104_18_ = ~(n_233 & ~(n_230 & in1_103_18_));
 assign in1_104_5_ = ~(n_238 & ~(n_230 & in1_103_5_));
 assign in1_104_2_ = ~(n_241 & n_236);
 assign in1_104_12_ = ~(n_231 & ~(n_230 & in1_103_12_));
 assign in1_104_1_ = ~(n_232 & ~(in1_101_0_ & in1_103_24_));
 assign in1_104_0_ = ~(n_235 & ~(n_230 & in1_103_0_));
 assign in1_104_11_ = ~(n_258 & n_237);
 assign n_259 = ~(in1_101_5_ & in1_103_24_);
 assign n_258 = ~(n_230 & in1_103_11_);
 assign n_257 = ~(in1_101_21_ & in1_103_24_);
 assign n_256 = ~(in1_101_16_ & in1_103_24_);
 assign n_255 = ~(in1_101_9_ & in1_103_24_);
 assign n_254 = ~(n_230 & in1_103_10_);
 assign n_253 = ~(in1_101_19_ & in1_103_24_);
 assign n_252 = ~(in1_101_8_ & in1_103_24_);
 assign n_251 = ~(in1_101_15_ & in1_103_24_);
 assign n_250 = ~(in1_101_14_ & in1_103_24_);
 assign n_249 = ~(in1_101_7_ & in1_103_24_);
 assign n_248 = ~(in1_101_6_ & in1_103_24_);
 assign n_247 = ~(n_230 & in1_103_7_);
 assign n_246 = ~(in1_101_22_ & in1_103_24_);
 assign n_245 = ~(in1_101_20_ & in1_103_24_);
 assign n_244 = ~(in1_101_18_ & in1_103_24_);
 assign n_243 = ~(in1_101_13_ & in1_103_24_);
 assign n_242 = ~(in1_101_3_ & in1_103_24_);
 assign n_241 = ~(n_230 & in1_103_2_);
 assign n_240 = ~(n_230 & in1_103_3_);
 assign n_239 = ~(in1_101_12_ & in1_103_24_);
 assign n_238 = ~(in1_101_4_ & in1_103_24_);
 assign n_237 = ~(in1_101_10_ & in1_103_24_);
 assign n_236 = ~(in1_101_1_ & in1_103_24_);
 assign n_235 = ~(in1_103_24_ & n_1548);
 assign n_234 = ~(in1_103_21_ & ~in1_103_24_);
 assign n_233 = ~(in1_101_17_ & in1_103_24_);
 assign n_232 = ~(n_230 & in1_103_1_);
 assign n_231 = ~(in1_101_11_ & in1_103_24_);
 assign n_230 = ~in1_103_24_;
 assign in1_107_8_ = ~(n_220 & ~(n_203 & in1_106_8_));
 assign in1_107_20_ = ~(n_224 & ~(n_203 & in1_106_20_));
 assign in1_107_17_ = ~(n_226 & ~(n_203 & in1_106_17_));
 assign in1_107_10_ = ~(n_225 & ~(n_203 & in1_106_10_));
 assign in1_107_16_ = ~(n_222 & ~(n_203 & in1_106_16_));
 assign in1_107_9_ = ~(n_223 & ~(n_203 & in1_106_9_));
 assign in1_107_23_ = ~(n_229 & ~(n_203 & in1_106_23_));
 assign in1_107_19_ = ~(n_216 & ~(n_203 & in1_106_19_));
 assign in1_107_15_ = ~(n_221 & ~(n_203 & in1_106_15_));
 assign in1_107_7_ = ~(n_219 & ~(in1_104_6_ & in1_106_24_));
 assign in1_107_6_ = ~(n_218 & ~(n_203 & in1_106_6_));
 assign in1_107_14_ = ~(n_213 & ~(in1_104_13_ & in1_106_24_));
 assign in1_107_13_ = ~(n_209 & ~(in1_104_12_ & in1_106_24_));
 assign in1_107_22_ = ~(n_227 & ~(n_203 & in1_106_22_));
 assign in1_107_21_ = ~(n_211 & ~(n_203 & in1_106_21_));
 assign in1_107_4_ = ~(n_215 & ~(n_203 & in1_106_4_));
 assign in1_107_3_ = ~(n_212 & ~(in1_104_2_ & in1_106_24_));
 assign in1_107_18_ = ~(n_207 & ~(n_203 & in1_106_18_));
 assign in1_107_5_ = ~(n_217 & ~(n_203 & in1_106_5_));
 assign in1_107_2_ = ~(n_214 & n_210);
 assign in1_107_12_ = ~(n_205 & ~(n_203 & in1_106_12_));
 assign in1_107_1_ = ~(n_206 & ~(in1_104_0_ & in1_106_24_));
 assign in1_107_0_ = ~(n_204 & n_208);
 assign in1_107_11_ = ~(n_228 & ~(in1_104_10_ & in1_106_24_));
 assign n_229 = ~(in1_104_22_ & in1_106_24_);
 assign n_228 = ~(n_203 & in1_106_11_);
 assign n_227 = ~(in1_104_21_ & in1_106_24_);
 assign n_226 = ~(in1_104_16_ & in1_106_24_);
 assign n_225 = ~(in1_104_9_ & in1_106_24_);
 assign n_224 = ~(in1_104_19_ & in1_106_24_);
 assign n_223 = ~(in1_104_8_ & in1_106_24_);
 assign n_222 = ~(in1_104_15_ & in1_106_24_);
 assign n_221 = ~(in1_104_14_ & in1_106_24_);
 assign n_220 = ~(in1_104_7_ & in1_106_24_);
 assign n_219 = ~(n_203 & in1_106_7_);
 assign n_218 = ~(in1_104_5_ & in1_106_24_);
 assign n_217 = ~(in1_104_4_ & in1_106_24_);
 assign n_216 = ~(in1_104_18_ & in1_106_24_);
 assign n_215 = ~(in1_104_3_ & in1_106_24_);
 assign n_214 = ~(n_203 & in1_106_2_);
 assign n_213 = ~(n_203 & in1_106_14_);
 assign n_212 = ~(n_203 & in1_106_3_);
 assign n_211 = ~(in1_104_20_ & in1_106_24_);
 assign n_210 = ~(in1_104_1_ & in1_106_24_);
 assign n_209 = ~(n_203 & in1_106_13_);
 assign n_208 = ~(in1_106_24_ & n_1537);
 assign n_207 = ~(in1_104_17_ & in1_106_24_);
 assign n_206 = ~(n_203 & in1_106_1_);
 assign n_205 = ~(in1_104_11_ & in1_106_24_);
 assign n_204 = ~(n_203 & in1_106_0_);
 assign n_203 = ~in1_106_24_;
 assign in1_110_8_ = ~(n_194 & ~(n_178 & n_1426));
 assign in1_110_20_ = ~(n_198 & ~(n_178 & in1_109_20_));
 assign in1_110_17_ = ~(n_200 & ~(n_178 & in1_109_17_));
 assign in1_110_10_ = ~(n_199 & ~(n_178 & n_1429));
 assign in1_110_16_ = ~(n_202 & ~(n_178 & in1_109_16_));
 assign in1_110_9_ = ~(n_197 & ~(n_178 & n_1452));
 assign in1_110_23_ = ~(n_196 & ~(n_178 & in1_109_23_));
 assign in1_110_19_ = ~(n_184 & ~(n_178 & in1_109_19_));
 assign in1_110_15_ = ~(n_195 & ~(n_178 & in1_109_15_));
 assign in1_110_7_ = ~(n_193 & ~(n_1455 & in1_109_24_));
 assign in1_110_6_ = ~(n_192 & ~(n_178 & n_1427));
 assign in1_110_14_ = ~(n_189 & ~(n_178 & in1_109_14_));
 assign in1_110_13_ = ~(n_187 & ~(n_178 & n_1412));
 assign in1_110_22_ = ~(n_201 & ~(n_178 & in1_109_22_));
 assign in1_110_21_ = ~(n_186 & ~(n_178 & in1_109_21_));
 assign in1_110_4_ = ~(n_188 & ~(n_178 & n_1432));
 assign in1_110_3_ = ~(n_183 & ~(n_178 & n_1434));
 assign in1_110_18_ = ~(n_182 & ~(n_178 & in1_109_18_));
 assign in1_110_5_ = ~(n_191 & ~(n_178 & n_1428));
 assign in1_110_2_ = ~(n_190 & ~(n_178 & n_1449));
 assign in1_110_12_ = ~(n_180 & ~(n_178 & n_1416));
 assign in1_110_1_ = ~(n_181 & ~(n_1467 & in1_109_24_));
 assign in1_110_0_ = ~(n_179 & ~(in1_109_24_ & n_1539));
 assign in1_110_11_ = ~(n_185 & ~(n_178 & n_1430));
 assign n_202 = ~(n_1421 & in1_109_24_);
 assign n_201 = ~(n_1442 & in1_109_24_);
 assign n_200 = ~(n_1456 & in1_109_24_);
 assign n_199 = ~(n_1443 & in1_109_24_);
 assign n_198 = ~(n_1450 & in1_109_24_);
 assign n_197 = ~(n_1451 & in1_109_24_);
 assign n_196 = ~(n_1439 & in1_109_24_);
 assign n_195 = ~(n_1422 & in1_109_24_);
 assign n_194 = ~(n_1409 & in1_109_24_);
 assign n_193 = ~(n_178 & n_1454);
 assign n_192 = ~(n_1410 & in1_109_24_);
 assign n_191 = ~(n_1425 & in1_109_24_);
 assign n_190 = ~(n_1448 & in1_109_24_);
 assign n_189 = ~(n_1436 & in1_109_24_);
 assign n_188 = ~(n_1431 & in1_109_24_);
 assign n_187 = ~(n_1435 & in1_109_24_);
 assign n_186 = ~(n_1444 & in1_109_24_);
 assign n_185 = ~(n_1420 & in1_109_24_);
 assign n_184 = ~(n_1441 & in1_109_24_);
 assign n_183 = ~(n_1433 & in1_109_24_);
 assign n_182 = ~(n_1445 & in1_109_24_);
 assign n_181 = ~(n_178 & in1_109_1_);
 assign n_180 = ~(n_1411 & in1_109_24_);
 assign n_179 = ~(n_178 & in1_109_0_);
 assign n_178 = ~in1_109_24_;
 assign in1_113_8_ = ~(n_169 & ~(n_150 & in1_112_8_));
 assign in1_113_20_ = ~(n_173 & ~(n_150 & in1_112_20_));
 assign in1_113_17_ = ~(n_175 & ~(n_150 & in1_112_17_));
 assign in1_113_10_ = ~(n_174 & ~(n_150 & in1_112_10_));
 assign in1_113_16_ = ~(n_171 & ~(n_150 & in1_112_16_));
 assign in1_113_9_ = ~(n_172 & ~(n_150 & in1_112_9_));
 assign in1_113_23_ = ~(n_177 & ~(n_150 & in1_112_23_));
 assign in1_113_19_ = ~(n_151 & ~(n_150 & in1_112_19_));
 assign in1_113_15_ = ~(n_170 & ~(n_150 & in1_112_15_));
 assign in1_113_7_ = ~(n_168 & ~(n_150 & in1_112_7_));
 assign in1_113_6_ = ~(n_166 & n_167);
 assign in1_113_14_ = ~(n_163 & ~(n_150 & in1_112_14_));
 assign in1_113_13_ = ~(n_157 & n_161);
 assign in1_113_22_ = ~(n_176 & ~(n_150 & in1_112_22_));
 assign in1_113_21_ = ~(n_160 & ~(n_150 & in1_112_21_));
 assign in1_113_4_ = ~(n_162 & ~(n_150 & in1_112_4_));
 assign in1_113_3_ = ~(n_156 & ~(n_150 & in1_112_3_));
 assign in1_113_18_ = ~(n_154 & ~(n_150 & in1_112_18_));
 assign in1_113_5_ = ~(n_165 & ~(n_150 & in1_112_5_));
 assign in1_113_2_ = ~(n_158 & ~(n_150 & in1_112_2_));
 assign in1_113_12_ = ~(n_152 & ~(n_150 & in1_112_12_));
 assign in1_113_1_ = ~(n_153 & ~(in1_110_0_ & in1_112_24_));
 assign in1_113_0_ = ~(n_164 & n_155);
 assign in1_113_11_ = ~(n_159 & ~(n_150 & in1_112_11_));
 assign n_177 = ~(in1_110_22_ & in1_112_24_);
 assign n_176 = ~(in1_110_21_ & in1_112_24_);
 assign n_175 = ~(in1_110_16_ & in1_112_24_);
 assign n_174 = ~(in1_110_9_ & in1_112_24_);
 assign n_173 = ~(in1_110_19_ & in1_112_24_);
 assign n_172 = ~(in1_110_8_ & in1_112_24_);
 assign n_171 = ~(in1_110_15_ & in1_112_24_);
 assign n_170 = ~(in1_110_14_ & in1_112_24_);
 assign n_169 = ~(in1_110_7_ & in1_112_24_);
 assign n_168 = ~(in1_110_6_ & in1_112_24_);
 assign n_167 = ~(in1_110_5_ & in1_112_24_);
 assign n_166 = ~(n_150 & in1_112_6_);
 assign n_165 = ~(in1_110_4_ & in1_112_24_);
 assign n_164 = ~(n_150 & in1_112_0_);
 assign n_163 = ~(in1_110_13_ & in1_112_24_);
 assign n_162 = ~(in1_110_3_ & in1_112_24_);
 assign n_161 = ~(in1_110_12_ & in1_112_24_);
 assign n_160 = ~(in1_110_20_ & in1_112_24_);
 assign n_159 = ~(in1_110_10_ & in1_112_24_);
 assign n_158 = ~(in1_110_1_ & in1_112_24_);
 assign n_157 = ~(n_150 & in1_112_13_);
 assign n_156 = ~(in1_110_2_ & in1_112_24_);
 assign n_155 = ~(in1_112_24_ & n_1523);
 assign n_154 = ~(in1_110_17_ & in1_112_24_);
 assign n_153 = ~(n_150 & in1_112_1_);
 assign n_152 = ~(in1_110_11_ & in1_112_24_);
 assign n_151 = ~(in1_110_18_ & in1_112_24_);
 assign n_150 = ~in1_112_24_;
 assign in1_116_8_ = ~(n_141 & ~(n_122 & in1_115_8_));
 assign in1_116_20_ = ~(n_145 & ~(n_122 & in1_115_20_));
 assign in1_116_17_ = ~(n_147 & ~(n_122 & in1_115_17_));
 assign in1_116_10_ = ~(n_146 & ~(in1_113_9_ & in1_115_24_));
 assign in1_116_16_ = ~(n_149 & ~(n_122 & in1_115_16_));
 assign in1_116_9_ = ~(n_144 & ~(in1_113_8_ & in1_115_24_));
 assign in1_116_23_ = ~(n_143 & ~(n_122 & in1_115_23_));
 assign in1_116_19_ = ~(n_137 & ~(n_122 & in1_115_19_));
 assign in1_116_15_ = ~(n_142 & ~(n_122 & in1_115_15_));
 assign in1_116_7_ = ~(n_140 & (in1_115_24_ | n_124));
 assign in1_116_6_ = ~(n_139 & ~(n_122 & in1_115_6_));
 assign in1_116_14_ = ~(n_136 & ~(n_122 & in1_115_14_));
 assign in1_116_13_ = ~(n_131 & ~(in1_113_12_ & in1_115_24_));
 assign in1_116_22_ = ~(n_148 & ~(n_122 & in1_115_22_));
 assign in1_116_21_ = ~(n_134 & ~(n_122 & in1_115_21_));
 assign in1_116_4_ = ~(n_135 & ~(n_122 & in1_115_4_));
 assign in1_116_3_ = ~(n_130 & ~(n_122 & in1_115_3_));
 assign in1_116_18_ = ~(n_128 & ~(n_122 & in1_115_18_));
 assign in1_116_5_ = ~(n_138 & ~(n_122 & in1_115_5_));
 assign in1_116_2_ = ~(n_132 & ~(n_122 & in1_115_2_));
 assign in1_116_12_ = ~(n_126 & ~(n_122 & in1_115_12_));
 assign in1_116_1_ = ~(n_127 & ~(in1_113_0_ & in1_115_24_));
 assign in1_116_0_ = ~(n_125 & n_129);
 assign in1_116_11_ = ~(n_133 & (in1_115_24_ | n_123));
 assign n_149 = ~(in1_113_15_ & in1_115_24_);
 assign n_148 = ~(in1_113_21_ & in1_115_24_);
 assign n_147 = ~(in1_113_16_ & in1_115_24_);
 assign n_146 = ~(n_122 & in1_115_10_);
 assign n_145 = ~(in1_113_19_ & in1_115_24_);
 assign n_144 = ~(n_122 & in1_115_9_);
 assign n_143 = ~(in1_113_22_ & in1_115_24_);
 assign n_142 = ~(in1_113_14_ & in1_115_24_);
 assign n_141 = ~(in1_113_7_ & in1_115_24_);
 assign n_140 = ~(in1_113_6_ & in1_115_24_);
 assign n_139 = ~(in1_113_5_ & in1_115_24_);
 assign n_138 = ~(in1_113_4_ & in1_115_24_);
 assign n_137 = ~(in1_113_18_ & in1_115_24_);
 assign n_136 = ~(in1_113_13_ & in1_115_24_);
 assign n_135 = ~(in1_113_3_ & in1_115_24_);
 assign n_134 = ~(in1_113_20_ & in1_115_24_);
 assign n_133 = ~(in1_113_10_ & in1_115_24_);
 assign n_132 = ~(in1_113_1_ & in1_115_24_);
 assign n_131 = ~(n_122 & in1_115_13_);
 assign n_130 = ~(in1_113_2_ & in1_115_24_);
 assign n_129 = ~(in1_115_24_ & n_1510);
 assign n_128 = ~(in1_113_17_ & in1_115_24_);
 assign n_127 = ~(n_122 & in1_115_1_);
 assign n_126 = ~(in1_113_11_ & in1_115_24_);
 assign n_125 = ~(n_122 & in1_115_0_);
 assign n_124 = ~in1_115_7_;
 assign n_123 = ~in1_115_11_;
 assign n_122 = ~in1_115_24_;
 assign in1_119_8_ = ~(n_111 & ~(n_95 & in1_118_8_));
 assign in1_119_20_ = ~(n_116 & ~(n_95 & in1_118_20_));
 assign in1_119_17_ = ~(n_119 & ~(n_95 & in1_118_17_));
 assign in1_119_10_ = ~(n_117 & ~(n_95 & in1_118_10_));
 assign in1_119_16_ = ~(n_113 & ~(n_95 & in1_118_16_));
 assign in1_119_9_ = ~(n_114 & n_115);
 assign in1_119_23_ = ~(n_121 & ~(n_95 & in1_118_23_));
 assign in1_119_19_ = ~(n_107 & ~(n_95 & in1_118_19_));
 assign in1_119_15_ = ~(n_112 & ~(n_95 & in1_118_15_));
 assign in1_119_7_ = ~(n_109 & n_110);
 assign in1_119_6_ = ~(n_108 & ~(n_95 & in1_118_6_));
 assign in1_119_14_ = ~(n_106 & ~(n_95 & in1_118_14_));
 assign in1_119_13_ = ~(n_102 & ~(n_95 & in1_118_13_));
 assign in1_119_22_ = ~(n_120 & ~(n_95 & in1_118_22_));
 assign in1_119_21_ = ~(n_101 & ~(n_95 & in1_118_21_));
 assign in1_119_4_ = ~(n_104 & ~(in1_116_3_ & in1_118_24_));
 assign in1_119_3_ = ~(n_103 & ~(in1_116_2_ & in1_118_24_));
 assign in1_119_18_ = ~(n_98 & ~(n_95 & in1_118_18_));
 assign in1_119_5_ = ~(n_118 & ~(in1_116_4_ & in1_118_24_));
 assign in1_119_2_ = ~(n_105 & ~(in1_116_1_ & in1_118_24_));
 assign in1_119_12_ = ~(n_96 & ~(n_95 & in1_118_12_));
 assign in1_119_1_ = ~(n_97 & ~(in1_116_0_ & in1_118_24_));
 assign in1_119_0_ = ~(n_99 & (in1_118_24_ | n_94));
 assign in1_119_11_ = ~(n_100 & ~(n_95 & in1_118_11_));
 assign n_121 = ~(in1_116_22_ & in1_118_24_);
 assign n_120 = ~(in1_116_21_ & in1_118_24_);
 assign n_119 = ~(in1_116_16_ & in1_118_24_);
 assign n_118 = ~(n_95 & in1_118_5_);
 assign n_117 = ~(in1_116_9_ & in1_118_24_);
 assign n_116 = ~(in1_116_19_ & in1_118_24_);
 assign n_115 = ~(in1_116_8_ & in1_118_24_);
 assign n_114 = ~(n_95 & in1_118_9_);
 assign n_113 = ~(in1_116_15_ & in1_118_24_);
 assign n_112 = ~(in1_116_14_ & in1_118_24_);
 assign n_111 = ~(in1_116_7_ & in1_118_24_);
 assign n_110 = ~(in1_116_6_ & in1_118_24_);
 assign n_109 = ~(n_95 & in1_118_7_);
 assign n_108 = ~(in1_116_5_ & in1_118_24_);
 assign n_107 = ~(in1_116_18_ & in1_118_24_);
 assign n_106 = ~(in1_116_13_ & in1_118_24_);
 assign n_105 = ~(n_95 & in1_118_2_);
 assign n_104 = ~(n_95 & in1_118_4_);
 assign n_103 = ~(n_95 & in1_118_3_);
 assign n_102 = ~(in1_116_12_ & in1_118_24_);
 assign n_101 = ~(in1_116_20_ & in1_118_24_);
 assign n_100 = ~(in1_116_10_ & in1_118_24_);
 assign n_99 = ~(in1_118_24_ & n_1547);
 assign n_98 = ~(in1_116_17_ & in1_118_24_);
 assign n_97 = ~(n_95 & in1_118_1_);
 assign n_96 = ~(in1_116_11_ & in1_118_24_);
 assign n_95 = ~in1_118_24_;
 assign n_94 = ~in1_118_0_;
 assign in1_122_8_ = ~(n_82 & ~(n_63 & in1_121_8_));
 assign in1_122_20_ = ~(n_87 & ~(n_63 & in1_121_20_));
 assign in1_122_17_ = ~(n_89 & n_91);
 assign in1_122_10_ = ~(n_88 & ~(n_63 & in1_121_10_));
 assign in1_122_16_ = ~(n_81 & n_84);
 assign in1_122_9_ = ~(n_85 & n_93);
 assign in1_122_23_ = ~(n_86 & ~(n_63 & in1_121_23_));
 assign in1_122_19_ = ~(n_76 & ~(n_63 & in1_121_19_));
 assign in1_122_15_ = ~(n_79 & n_83);
 assign in1_122_7_ = ~(n_80 & ~(n_63 & in1_121_7_));
 assign in1_122_6_ = ~(n_71 & ~(n_63 & in1_121_6_));
 assign in1_122_14_ = ~(n_75 & ~(n_63 & in1_121_14_));
 assign in1_122_13_ = ~(n_72 & ~(n_63 & in1_121_13_));
 assign in1_122_22_ = ~(n_92 & ~(n_63 & in1_121_22_));
 assign in1_122_21_ = ~(n_78 & ~(n_63 & in1_121_21_));
 assign in1_122_4_ = ~(n_74 & ~(n_63 & in1_121_4_));
 assign in1_122_3_ = ~(n_68 & ~(n_63 & in1_121_3_));
 assign in1_122_18_ = ~(n_67 & ~(n_63 & in1_121_18_));
 assign in1_122_5_ = ~(n_90 & n_77);
 assign in1_122_2_ = ~(n_73 & n_69);
 assign in1_122_12_ = ~(n_65 & ~(n_63 & in1_121_12_));
 assign in1_122_1_ = ~(n_66 & ~(in1_119_0_ & in1_121_24_));
 assign in1_122_0_ = ~(n_64 & ~(in1_121_24_ & n_1402));
 assign in1_122_11_ = ~(n_70 & ~(n_63 & in1_121_11_));
 assign n_93 = ~(in1_119_8_ & in1_121_24_);
 assign n_92 = ~(in1_119_21_ & in1_121_24_);
 assign n_91 = ~(in1_119_16_ & in1_121_24_);
 assign n_90 = ~(n_63 & in1_121_5_);
 assign n_89 = ~(n_63 & in1_121_17_);
 assign n_88 = ~(in1_119_9_ & in1_121_24_);
 assign n_87 = ~(in1_119_19_ & in1_121_24_);
 assign n_86 = ~(in1_119_22_ & in1_121_24_);
 assign n_85 = ~(n_63 & in1_121_9_);
 assign n_84 = ~(in1_119_15_ & in1_121_24_);
 assign n_83 = ~(in1_119_14_ & in1_121_24_);
 assign n_82 = ~(in1_119_7_ & in1_121_24_);
 assign n_81 = ~(n_63 & in1_121_16_);
 assign n_80 = ~(in1_119_6_ & in1_121_24_);
 assign n_79 = ~(n_63 & in1_121_15_);
 assign n_78 = ~(in1_119_20_ & in1_121_24_);
 assign n_77 = ~(in1_119_4_ & in1_121_24_);
 assign n_76 = ~(in1_119_18_ & in1_121_24_);
 assign n_75 = ~(in1_119_13_ & in1_121_24_);
 assign n_74 = ~(in1_119_3_ & in1_121_24_);
 assign n_73 = ~(n_63 & in1_121_2_);
 assign n_72 = ~(in1_119_12_ & in1_121_24_);
 assign n_71 = ~(in1_119_5_ & in1_121_24_);
 assign n_70 = ~(in1_119_10_ & in1_121_24_);
 assign n_69 = ~(in1_119_1_ & in1_121_24_);
 assign n_68 = ~(in1_119_2_ & in1_121_24_);
 assign n_67 = ~(in1_119_17_ & in1_121_24_);
 assign n_66 = ~(n_63 & in1_121_1_);
 assign n_65 = ~(in1_119_11_ & in1_121_24_);
 assign n_64 = ~(n_63 & in1_121_0_);
 assign n_63 = ~in1_121_24_;
 assign in1_125_8_ = ~(n_52 & ~(n_35 & in1_124_8_));
 assign in1_125_20_ = ~(n_57 & ~(n_35 & in1_124_20_));
 assign in1_125_17_ = ~(n_59 & ~(n_35 & in1_124_17_));
 assign in1_125_10_ = ~(n_58 & ~(n_35 & in1_124_10_));
 assign in1_125_16_ = ~(n_51 & n_54);
 assign in1_125_9_ = ~(n_55 & n_56);
 assign in1_125_23_ = ~(n_62 & ~(n_35 & in1_124_23_));
 assign in1_125_19_ = ~(n_47 & ~(n_35 & in1_124_19_));
 assign in1_125_15_ = ~(n_53 & ~(n_35 & in1_124_15_));
 assign in1_125_7_ = ~(n_50 & ~(in1_122_6_ & in1_124_24_));
 assign in1_125_6_ = ~(n_36 & ~(n_35 & in1_124_6_));
 assign in1_125_14_ = ~(n_46 & ~(n_35 & in1_124_14_));
 assign in1_125_13_ = ~(n_41 & ~(in1_122_12_ & in1_124_24_));
 assign in1_125_22_ = ~(n_60 & ~(n_35 & in1_124_22_));
 assign in1_125_21_ = ~(n_43 & ~(n_35 & in1_124_21_));
 assign in1_125_4_ = ~(n_45 & ~(n_35 & in1_124_4_));
 assign in1_125_3_ = ~(n_40 & ~(n_35 & in1_124_3_));
 assign in1_125_18_ = ~(n_39 & ~(n_35 & in1_124_18_));
 assign in1_125_5_ = ~(n_48 & ~(n_35 & in1_124_5_));
 assign in1_125_2_ = ~(n_44 & n_42);
 assign in1_125_12_ = ~(n_37 & ~(n_35 & in1_124_12_));
 assign in1_125_1_ = ~(n_38 & ~(in1_122_0_ & in1_124_24_));
 assign in1_125_0_ = ~(n_49 & ~(in1_124_24_ & n_1598));
 assign in1_125_11_ = ~(n_61 & ~(in1_122_10_ & in1_124_24_));
 assign n_62 = ~(in1_122_22_ & in1_124_24_);
 assign n_61 = ~(n_35 & in1_124_11_);
 assign n_60 = ~(in1_122_21_ & in1_124_24_);
 assign n_59 = ~(in1_122_16_ & in1_124_24_);
 assign n_58 = ~(in1_122_9_ & in1_124_24_);
 assign n_57 = ~(in1_122_19_ & in1_124_24_);
 assign n_56 = ~(in1_122_8_ & in1_124_24_);
 assign n_55 = ~(n_35 & in1_124_9_);
 assign n_54 = ~(in1_122_15_ & in1_124_24_);
 assign n_53 = ~(in1_122_14_ & in1_124_24_);
 assign n_52 = ~(in1_122_7_ & in1_124_24_);
 assign n_51 = ~(n_35 & in1_124_16_);
 assign n_50 = ~(n_35 & in1_124_7_);
 assign n_49 = ~(n_35 & in1_124_0_);
 assign n_48 = ~(in1_122_4_ & in1_124_24_);
 assign n_47 = ~(in1_122_18_ & in1_124_24_);
 assign n_46 = ~(in1_122_13_ & in1_124_24_);
 assign n_45 = ~(in1_122_3_ & in1_124_24_);
 assign n_44 = ~(n_35 & in1_124_2_);
 assign n_43 = ~(in1_122_20_ & in1_124_24_);
 assign n_42 = ~(in1_122_1_ & in1_124_24_);
 assign n_41 = ~(n_35 & in1_124_13_);
 assign n_40 = ~(in1_122_2_ & in1_124_24_);
 assign n_39 = ~(in1_122_17_ & in1_124_24_);
 assign n_38 = ~(n_35 & in1_124_1_);
 assign n_37 = ~(in1_122_11_ & in1_124_24_);
 assign n_36 = ~(in1_122_5_ & in1_124_24_);
 assign n_35 = ~in1_124_24_;
 assign in1_128_8_ = ~(n_26 & ~(n_9 & in1_127_8_));
 assign in1_128_20_ = ~(n_30 & ~(n_9 & in1_127_20_));
 assign in1_128_17_ = ~(n_33 & ~(n_9 & in1_127_17_));
 assign in1_128_10_ = ~(n_31 & ~(n_9 & in1_127_10_));
 assign in1_128_16_ = ~(n_34 & ~(n_9 & in1_127_16_));
 assign in1_128_9_ = ~(n_29 & ~(n_9 & in1_127_9_));
 assign in1_128_23_ = ((in1_127_23_ & ~in1_127_24_) | (in1_125_22_ & in1_127_24_));
 assign in1_128_19_ = ~(n_22 & ~(n_9 & in1_127_19_));
 assign in1_128_15_ = ~(n_27 & ~(n_9 & in1_127_15_));
 assign in1_128_7_ = ~(n_25 & ~(in1_125_6_ & in1_127_24_));
 assign in1_128_6_ = ~(n_24 & ~(n_9 & in1_127_6_));
 assign in1_128_14_ = ~(n_21 & ~(n_9 & in1_127_14_));
 assign in1_128_13_ = ~(n_14 & n_18);
 assign in1_128_22_ = ~(n_28 & ~(n_9 & in1_127_22_));
 assign in1_128_21_ = ~(n_17 & ~(n_9 & in1_127_21_));
 assign in1_128_4_ = ~(n_20 & ~(n_9 & in1_127_4_));
 assign in1_128_3_ = ~(n_19 & ~(in1_125_2_ & in1_127_24_));
 assign in1_128_18_ = ~(n_12 & ~(n_9 & in1_127_18_));
 assign in1_128_5_ = ~(n_32 & n_23);
 assign in1_128_2_ = ~(n_15 & ~(n_9 & in1_127_2_));
 assign in1_128_12_ = ~(n_10 & ~(n_9 & in1_127_12_));
 assign in1_128_1_ = ~(n_11 & ~(in1_125_0_ & in1_127_24_));
 assign in1_128_0_ = ~(n_13 & (in1_127_24_ | n_8));
 assign in1_128_11_ = ~(n_16 & ~(n_9 & in1_127_11_));
 assign n_34 = ~(in1_125_15_ & in1_127_24_);
 assign n_33 = ~(in1_125_16_ & in1_127_24_);
 assign n_32 = ~(n_9 & in1_127_5_);
 assign n_31 = ~(in1_125_9_ & in1_127_24_);
 assign n_30 = ~(in1_125_19_ & in1_127_24_);
 assign n_29 = ~(in1_125_8_ & in1_127_24_);
 assign n_28 = ~(in1_125_21_ & in1_127_24_);
 assign n_27 = ~(in1_125_14_ & in1_127_24_);
 assign n_26 = ~(in1_125_7_ & in1_127_24_);
 assign n_25 = ~(n_9 & in1_127_7_);
 assign n_24 = ~(in1_125_5_ & in1_127_24_);
 assign n_23 = ~(in1_125_4_ & in1_127_24_);
 assign n_22 = ~(in1_125_18_ & in1_127_24_);
 assign n_21 = ~(in1_125_13_ & in1_127_24_);
 assign n_20 = ~(in1_125_3_ & in1_127_24_);
 assign n_19 = ~(n_9 & in1_127_3_);
 assign n_18 = ~(in1_125_12_ & in1_127_24_);
 assign n_17 = ~(in1_125_20_ & in1_127_24_);
 assign n_16 = ~(in1_125_10_ & in1_127_24_);
 assign n_15 = ~(in1_125_1_ & in1_127_24_);
 assign n_14 = ~(n_9 & in1_127_13_);
 assign n_13 = ~(in1_127_24_ & n_1576);
 assign n_12 = ~(in1_125_17_ & in1_127_24_);
 assign n_11 = ~(n_9 & in1_127_1_);
 assign n_10 = ~(in1_125_11_ & in1_127_24_);
 assign n_9 = ~in1_127_24_;
 assign n_8 = ~in1_127_0_;
 assign in1_131_8_ = ((in1_130_8_ & ~in1_130_24_) | (in1_128_7_ & in1_130_24_));
 assign in1_131_20_ = ((in1_130_20_ & ~in1_130_24_) | (in1_128_19_ & in1_130_24_));
 assign in1_131_17_ = ((in1_130_17_ & ~in1_130_24_) | (in1_128_16_ & in1_130_24_));
 assign in1_131_10_ = ((in1_130_10_ & ~in1_130_24_) | (in1_128_9_ & in1_130_24_));
 assign in1_131_16_ = ((in1_130_16_ & ~in1_130_24_) | (in1_128_15_ & in1_130_24_));
 assign in1_131_9_ = ((in1_130_9_ & ~in1_130_24_) | (in1_128_8_ & in1_130_24_));
 assign in1_131_23_ = ((in1_130_23_ & ~in1_130_24_) | (in1_128_22_ & in1_130_24_));
 assign in1_131_19_ = ~(n_5 & ~(n_1 & in1_130_19_));
 assign in1_131_15_ = ((in1_130_15_ & ~in1_130_24_) | (in1_128_14_ & in1_130_24_));
 assign in1_131_7_ = ((in1_130_7_ & ~in1_130_24_) | (in1_128_6_ & in1_130_24_));
 assign in1_131_6_ = ((in1_130_6_ & ~in1_130_24_) | (in1_128_5_ & in1_130_24_));
 assign in1_131_14_ = ((in1_130_14_ & ~in1_130_24_) | (in1_128_13_ & in1_130_24_));
 assign in1_131_13_ = ((in1_130_13_ & ~in1_130_24_) | (in1_128_12_ & in1_130_24_));
 assign in1_131_22_ = ~(n_7 & ~(n_1 & in1_130_22_));
 assign in1_131_21_ = ((in1_130_21_ & ~in1_130_24_) | (in1_128_20_ & in1_130_24_));
 assign in1_131_4_ = ~(n_4 & ~(n_1 & in1_130_4_));
 assign in1_131_3_ = ((in1_130_3_ & ~in1_130_24_) | (in1_128_2_ & in1_130_24_));
 assign in1_131_18_ = ((in1_130_18_ & ~in1_130_24_) | (in1_128_17_ & in1_130_24_));
 assign in1_131_5_ = ((in1_130_5_ & ~in1_130_24_) | (in1_128_4_ & in1_130_24_));
 assign in1_131_2_ = ~(n_3 & ~(n_1 & in1_130_2_));
 assign in1_131_12_ = ((in1_130_12_ & ~in1_130_24_) | (in1_128_11_ & in1_130_24_));
 assign in1_131_1_ = ~(n_6 & ~(n_1 & in1_130_1_));
 assign in1_131_0_ = ~(n_2 & (in1_130_24_ | n_0));
 assign in1_131_11_ = ((in1_130_11_ & ~in1_130_24_) | (in1_128_10_ & in1_130_24_));
 assign n_7 = ~(in1_128_21_ & in1_130_24_);
 assign n_6 = ~(in1_128_0_ & in1_130_24_);
 assign n_5 = ~(in1_128_18_ & in1_130_24_);
 assign n_4 = ~(in1_128_3_ & in1_130_24_);
 assign n_3 = ~(in1_128_1_ & in1_130_24_);
 assign n_2 = ~(in1_130_24_ & n_1574);
 assign n_1 = ~in1_130_24_;
 assign n_0 = ~in1_130_0_;
 assign in1_134_8_ = ((in1_133_8_ & ~in1_133_24_) | (in1_131_7_ & in1_133_24_));
 assign in1_134_20_ = ((in1_133_20_ & ~in1_133_24_) | (in1_131_19_ & in1_133_24_));
 assign in1_134_17_ = ((in1_133_17_ & ~in1_133_24_) | (in1_131_16_ & in1_133_24_));
 assign in1_134_10_ = ((in1_133_10_ & ~in1_133_24_) | (in1_131_9_ & in1_133_24_));
 assign in1_134_16_ = ((in1_133_16_ & ~in1_133_24_) | (in1_131_15_ & in1_133_24_));
 assign in1_134_9_ = ((in1_133_9_ & ~in1_133_24_) | (in1_131_8_ & in1_133_24_));
 assign in1_134_23_ = ((in1_133_23_ & ~in1_133_24_) | (in1_131_22_ & in1_133_24_));
 assign in1_134_19_ = ((in1_133_19_ & ~in1_133_24_) | (in1_131_18_ & in1_133_24_));
 assign in1_134_15_ = ((in1_133_15_ & ~in1_133_24_) | (in1_131_14_ & in1_133_24_));
 assign in1_134_7_ = ((in1_133_7_ & ~in1_133_24_) | (in1_131_6_ & in1_133_24_));
 assign in1_134_6_ = ((in1_133_6_ & ~in1_133_24_) | (in1_131_5_ & in1_133_24_));
 assign in1_134_14_ = ((in1_133_14_ & ~in1_133_24_) | (in1_131_13_ & in1_133_24_));
 assign in1_134_13_ = ((in1_133_13_ & ~in1_133_24_) | (in1_131_12_ & in1_133_24_));
 assign in1_134_22_ = ((in1_133_22_ & ~in1_133_24_) | (in1_131_21_ & in1_133_24_));
 assign in1_134_21_ = ((in1_133_21_ & ~in1_133_24_) | (in1_131_20_ & in1_133_24_));
 assign in1_134_4_ = ((in1_133_4_ & ~in1_133_24_) | (in1_131_3_ & in1_133_24_));
 assign in1_134_3_ = ((in1_133_3_ & ~in1_133_24_) | (in1_131_2_ & in1_133_24_));
 assign in1_134_18_ = ((in1_133_18_ & ~in1_133_24_) | (in1_131_17_ & in1_133_24_));
 assign in1_134_5_ = ((in1_133_5_ & ~in1_133_24_) | (in1_131_4_ & in1_133_24_));
 assign in1_134_2_ = ((in1_133_2_ & ~in1_133_24_) | (in1_131_1_ & in1_133_24_));
 assign in1_134_12_ = ((in1_133_12_ & ~in1_133_24_) | (in1_131_11_ & in1_133_24_));
 assign in1_134_1_ = ((in1_133_1_ & ~in1_133_24_) | (in1_131_0_ & in1_133_24_));
 assign in1_134_0_ = ((in1_133_0_ & ~in1_133_24_) | (n_1531 & in1_133_24_));
 assign in1_134_11_ = ((in1_133_11_ & ~in1_133_24_) | (in1_131_10_ & in1_133_24_));
 assign in1_137_8_ = ((in1_136_8_ & ~in1_136_24_) | (in1_134_7_ & in1_136_24_));
 assign in1_137_20_ = ((in1_136_20_ & ~in1_136_24_) | (in1_134_19_ & in1_136_24_));
 assign in1_137_17_ = ((in1_136_17_ & ~in1_136_24_) | (in1_134_16_ & in1_136_24_));
 assign in1_137_10_ = ((in1_136_10_ & ~in1_136_24_) | (in1_134_9_ & in1_136_24_));
 assign in1_137_16_ = ((in1_136_16_ & ~in1_136_24_) | (in1_134_15_ & in1_136_24_));
 assign in1_137_9_ = ((in1_136_9_ & ~in1_136_24_) | (in1_134_8_ & in1_136_24_));
 assign in1_137_23_ = ((in1_136_23_ & ~in1_136_24_) | (in1_134_22_ & in1_136_24_));
 assign in1_137_19_ = ((in1_136_19_ & ~in1_136_24_) | (in1_134_18_ & in1_136_24_));
 assign in1_137_15_ = ((in1_136_15_ & ~in1_136_24_) | (in1_134_14_ & in1_136_24_));
 assign in1_137_7_ = ((in1_136_7_ & ~in1_136_24_) | (in1_134_6_ & in1_136_24_));
 assign in1_137_6_ = ((in1_136_6_ & ~in1_136_24_) | (in1_134_5_ & in1_136_24_));
 assign in1_137_14_ = ((in1_136_14_ & ~in1_136_24_) | (in1_134_13_ & in1_136_24_));
 assign in1_137_13_ = ((in1_136_13_ & ~in1_136_24_) | (in1_134_12_ & in1_136_24_));
 assign in1_137_22_ = ((in1_136_22_ & ~in1_136_24_) | (in1_134_21_ & in1_136_24_));
 assign in1_137_21_ = ((in1_136_21_ & ~in1_136_24_) | (in1_134_20_ & in1_136_24_));
 assign in1_137_4_ = ((in1_136_4_ & ~in1_136_24_) | (in1_134_3_ & in1_136_24_));
 assign in1_137_3_ = ((in1_136_3_ & ~in1_136_24_) | (in1_134_2_ & in1_136_24_));
 assign in1_137_18_ = ((in1_136_18_ & ~in1_136_24_) | (in1_134_17_ & in1_136_24_));
 assign in1_137_5_ = ((in1_136_5_ & ~in1_136_24_) | (in1_134_4_ & in1_136_24_));
 assign in1_137_2_ = ((in1_136_2_ & ~in1_136_24_) | (in1_134_1_ & in1_136_24_));
 assign in1_137_12_ = ((in1_136_12_ & ~in1_136_24_) | (in1_134_11_ & in1_136_24_));
 assign in1_137_1_ = ((in1_136_1_ & ~in1_136_24_) | (in1_134_0_ & in1_136_24_));
 assign in1_137_0_ = ((in1_136_0_ & ~in1_136_24_) | (n_1554 & in1_136_24_));
 assign in1_137_11_ = ((in1_136_11_ & ~in1_136_24_) | (in1_134_10_ & in1_136_24_));
 assign in1_140_8_ = ((in1_139_8_ & ~in1_139_24_) | (in1_137_7_ & in1_139_24_));
 assign in1_140_20_ = ((in1_139_20_ & ~in1_139_24_) | (in1_137_19_ & in1_139_24_));
 assign in1_140_17_ = ((in1_139_17_ & ~in1_139_24_) | (in1_137_16_ & in1_139_24_));
 assign in1_140_10_ = ((in1_139_10_ & ~in1_139_24_) | (in1_137_9_ & in1_139_24_));
 assign in1_140_16_ = ((in1_139_16_ & ~in1_139_24_) | (in1_137_15_ & in1_139_24_));
 assign in1_140_9_ = ((in1_139_9_ & ~in1_139_24_) | (in1_137_8_ & in1_139_24_));
 assign in1_140_23_ = ((in1_139_23_ & ~in1_139_24_) | (in1_137_22_ & in1_139_24_));
 assign in1_140_19_ = ((in1_139_19_ & ~in1_139_24_) | (in1_137_18_ & in1_139_24_));
 assign in1_140_15_ = ((in1_139_15_ & ~in1_139_24_) | (in1_137_14_ & in1_139_24_));
 assign in1_140_7_ = ((in1_139_7_ & ~in1_139_24_) | (in1_137_6_ & in1_139_24_));
 assign in1_140_6_ = ((in1_139_6_ & ~in1_139_24_) | (in1_137_5_ & in1_139_24_));
 assign in1_140_14_ = ((in1_139_14_ & ~in1_139_24_) | (in1_137_13_ & in1_139_24_));
 assign in1_140_13_ = ((in1_139_13_ & ~in1_139_24_) | (in1_137_12_ & in1_139_24_));
 assign in1_140_22_ = ((in1_139_22_ & ~in1_139_24_) | (in1_137_21_ & in1_139_24_));
 assign in1_140_21_ = ((in1_139_21_ & ~in1_139_24_) | (in1_137_20_ & in1_139_24_));
 assign in1_140_4_ = ((in1_139_4_ & ~in1_139_24_) | (in1_137_3_ & in1_139_24_));
 assign in1_140_3_ = ((in1_139_3_ & ~in1_139_24_) | (in1_137_2_ & in1_139_24_));
 assign in1_140_18_ = ((in1_139_18_ & ~in1_139_24_) | (in1_137_17_ & in1_139_24_));
 assign in1_140_5_ = ((in1_139_5_ & ~in1_139_24_) | (in1_137_4_ & in1_139_24_));
 assign in1_140_2_ = ((in1_139_2_ & ~in1_139_24_) | (in1_137_1_ & in1_139_24_));
 assign in1_140_12_ = ((in1_139_12_ & ~in1_139_24_) | (in1_137_11_ & in1_139_24_));
 assign in1_140_1_ = ((in1_139_1_ & ~in1_139_24_) | (in1_137_0_ & in1_139_24_));
 assign in1_140_0_ = ((in1_139_0_ & ~in1_139_24_) | (n_1471 & in1_139_24_));
 assign in1_140_11_ = ((in1_139_11_ & ~in1_139_24_) | (in1_137_10_ & in1_139_24_));
 assign in1_143_8_ = ((in1_142_8_ & ~in1_142_24_) | (in1_140_7_ & in1_142_24_));
 assign in1_143_20_ = ((in1_142_20_ & ~in1_142_24_) | (in1_140_19_ & in1_142_24_));
 assign in1_143_17_ = ((in1_142_17_ & ~in1_142_24_) | (in1_140_16_ & in1_142_24_));
 assign in1_143_10_ = ((in1_142_10_ & ~in1_142_24_) | (in1_140_9_ & in1_142_24_));
 assign in1_143_16_ = ((in1_142_16_ & ~in1_142_24_) | (in1_140_15_ & in1_142_24_));
 assign in1_143_9_ = ((in1_142_9_ & ~in1_142_24_) | (in1_140_8_ & in1_142_24_));
 assign in1_143_23_ = ((in1_142_23_ & ~in1_142_24_) | (in1_140_22_ & in1_142_24_));
 assign in1_143_19_ = ((in1_142_19_ & ~in1_142_24_) | (in1_140_18_ & in1_142_24_));
 assign in1_143_15_ = ((in1_142_15_ & ~in1_142_24_) | (in1_140_14_ & in1_142_24_));
 assign in1_143_7_ = ((in1_142_7_ & ~in1_142_24_) | (in1_140_6_ & in1_142_24_));
 assign in1_143_6_ = ((in1_142_6_ & ~in1_142_24_) | (in1_140_5_ & in1_142_24_));
 assign in1_143_14_ = ((in1_142_14_ & ~in1_142_24_) | (in1_140_13_ & in1_142_24_));
 assign in1_143_13_ = ((in1_142_13_ & ~in1_142_24_) | (in1_140_12_ & in1_142_24_));
 assign in1_143_22_ = ((in1_142_22_ & ~in1_142_24_) | (in1_140_21_ & in1_142_24_));
 assign in1_143_21_ = ((in1_142_21_ & ~in1_142_24_) | (in1_140_20_ & in1_142_24_));
 assign in1_143_4_ = ((in1_142_4_ & ~in1_142_24_) | (in1_140_3_ & in1_142_24_));
 assign in1_143_3_ = ((in1_142_3_ & ~in1_142_24_) | (in1_140_2_ & in1_142_24_));
 assign in1_143_18_ = ((in1_142_18_ & ~in1_142_24_) | (in1_140_17_ & in1_142_24_));
 assign in1_143_5_ = ((in1_142_5_ & ~in1_142_24_) | (in1_140_4_ & in1_142_24_));
 assign in1_143_2_ = ((in1_142_2_ & ~in1_142_24_) | (in1_140_1_ & in1_142_24_));
 assign in1_143_12_ = ((in1_142_12_ & ~in1_142_24_) | (in1_140_11_ & in1_142_24_));
 assign in1_143_1_ = ((in1_142_1_ & ~in1_142_24_) | (in1_140_0_ & in1_142_24_));
 assign in1_143_0_ = ((in1_142_0_ & ~in1_142_24_) | (n_1400 & in1_142_24_));
 assign in1_143_11_ = ((in1_142_11_ & ~in1_142_24_) | (in1_140_10_ & in1_142_24_));
 assign in1_1_24_ = ~(sub_217_2_n_25 & sub_217_2_n_2);
 assign sub_217_2_n_25 = ~(sub_217_2_n_23 | sub_217_2_n_21);
 assign sub_217_2_n_24 = ~(sub_217_2_n_22 & sub_217_2_n_12);
 assign sub_217_2_n_23 = ~(sub_217_2_n_17 & sub_217_2_n_19);
 assign sub_217_2_n_22 = ~(sub_217_2_n_16 | {in2[3]});
 assign sub_217_2_n_21 = ~(sub_217_2_n_15 & sub_217_2_n_18);
 assign in1_1_0_ = ~(sub_217_2_n_1 & sub_217_2_n_0);
 assign sub_217_2_n_19 = ~(sub_217_2_n_8 | sub_217_2_n_9);
 assign sub_217_2_n_18 = ~(sub_217_2_n_5 | sub_217_2_n_7);
 assign sub_217_2_n_17 = ~(sub_217_2_n_3 | sub_217_2_n_6);
 assign sub_217_2_n_16 = ~(sub_217_2_n_14 & sub_217_2_n_13);
 assign sub_217_2_n_15 = ~(sub_217_2_n_10 | sub_217_2_n_4);
 assign sub_217_2_n_14 = ~({in2[4]} | {in2[5]});
 assign sub_217_2_n_13 = ~({in2[14]} | {in2[15]});
 assign sub_217_2_n_12 = ~({in2[1]} | {in2[2]});
 assign sub_217_2_n_10 = ({in2[16]} | {in2[17]});
 assign sub_217_2_n_9 = ({in2[12]} | {in2[13]});
 assign sub_217_2_n_8 = ({in2[10]} | {in2[11]});
 assign sub_217_2_n_7 = ({in2[22]} | {in2[23]});
 assign sub_217_2_n_6 = ({in2[8]} | {in2[9]});
 assign sub_217_2_n_5 = ({in2[20]} | {in2[21]});
 assign sub_217_2_n_4 = ({in2[18]} | {in2[19]});
 assign sub_217_2_n_3 = ({in2[6]} | {in2[7]});
 assign sub_217_2_n_2 = ~(sub_217_2_n_24 | ~sub_217_2_n_0);
 assign sub_217_2_n_1 = ~({in1[48]} & ~{in2[0]});
 assign sub_217_2_n_0 = ~({in2[0]} & ~{in1[48]});
 assign in1_4_24_ = ~(sub_236_2_n_30 & (sub_236_2_n_27 | in1_2_0_));
 assign in1_4_1_ = ~((sub_236_2_n_29 & ~in1_2_0_) | (sub_236_2_n_28 & in1_2_0_));
 assign sub_236_2_n_30 = ~(sub_236_2_n_25 | (sub_236_2_n_23 | sub_236_2_n_26));
 assign sub_236_2_n_29 = ~sub_236_2_n_28;
 assign sub_236_2_n_28 = (sub_236_2_n_11 ^ sub_236_2_n_7);
 assign sub_236_2_n_27 = ~({in2[1]} | (sub_236_2_n_8 & {in2[0]}));
 assign sub_236_2_n_26 = ~(sub_236_2_n_11 | sub_236_2_n_7);
 assign sub_236_2_n_25 = ~(sub_236_2_n_24 & sub_236_2_n_22);
 assign sub_236_2_n_24 = ~(sub_236_2_n_17 | sub_236_2_n_18);
 assign sub_236_2_n_23 = ~(sub_236_2_n_19 & sub_236_2_n_16);
 assign sub_236_2_n_22 = ~(sub_236_2_n_20 | sub_236_2_n_1);
 assign in1_4_0_ = ~(sub_236_2_n_0 & sub_236_2_n_11);
 assign sub_236_2_n_20 = ~(sub_236_2_n_14 & sub_236_2_n_15);
 assign sub_236_2_n_19 = ~(sub_236_2_n_3 | sub_236_2_n_4);
 assign sub_236_2_n_18 = ~(sub_236_2_n_12 & sub_236_2_n_13);
 assign sub_236_2_n_17 = ~(sub_236_2_n_9 & sub_236_2_n_10);
 assign sub_236_2_n_16 = ~(sub_236_2_n_5 | sub_236_2_n_2);
 assign sub_236_2_n_15 = ~({in2[22]} | {in2[23]});
 assign sub_236_2_n_14 = ~({in2[20]} | {in2[21]});
 assign sub_236_2_n_13 = ~({in2[16]} | {in2[17]});
 assign sub_236_2_n_12 = ~({in2[14]} | {in2[15]});
 assign sub_236_2_n_10 = ~({in2[6]} | {in2[7]});
 assign sub_236_2_n_9 = ~({in2[4]} | {in2[5]});
 assign sub_236_2_n_11 = ~(sub_236_2_n_8 & {in2[0]});
 assign sub_236_2_n_8 = ~{in1[47]};
 assign sub_236_2_n_7 = ~{in2[1]};
 assign sub_236_2_n_5 = ({in2[12]} | {in2[13]});
 assign sub_236_2_n_4 = ({in2[8]} | {in2[9]});
 assign sub_236_2_n_3 = ({in2[2]} | {in2[3]});
 assign sub_236_2_n_2 = ({in2[18]} | {in2[19]});
 assign sub_236_2_n_1 = ({in2[10]} | {in2[11]});
 assign sub_236_2_n_0 = ~({in1[47]} & ~{in2[0]});
 assign in1_7_24_ = ~(sub_255_2_n_40 & (sub_255_2_n_39 | sub_255_2_n_28));
 assign in1_7_2_ = ~((sub_255_2_n_35 & ~sub_255_2_n_26) | (sub_255_2_n_41 & sub_255_2_n_26));
 assign sub_255_2_n_41 = ~sub_255_2_n_35;
 assign sub_255_2_n_40 = ~(sub_255_2_n_17 | ~sub_255_2_n_36);
 assign sub_255_2_n_39 = ~(sub_255_2_n_37 | ~sub_255_2_n_38);
 assign sub_255_2_n_38 = ~(sub_255_2_n_33 | {in2[3]});
 assign sub_255_2_n_37 = ~(in1_5_0_ | ~sub_255_2_n_32);
 assign sub_255_2_n_36 = ~(sub_255_2_n_31 | sub_255_2_n_30);
 assign sub_255_2_n_35 = ~(sub_255_2_n_3 | sub_255_2_n_0);
 assign in1_7_1_ = ~(in1_5_0_ ^ ({in2[1]} ^ sub_255_2_n_1));
 assign sub_255_2_n_33 = ~(sub_255_2_n_1 | ~{in2[1]});
 assign sub_255_2_n_32 = ~(sub_255_2_n_1 & ~{in2[1]});
 assign sub_255_2_n_31 = ~(sub_255_2_n_29 & sub_255_2_n_25);
 assign sub_255_2_n_30 = ~(sub_255_2_n_21 & sub_255_2_n_24);
 assign sub_255_2_n_29 = ~(sub_255_2_n_22 | sub_255_2_n_23);
 assign sub_255_2_n_28 = ~(sub_255_2_n_11 | ~sub_255_2_n_15);
 assign in1_7_0_ = ~(sub_255_2_n_2 & sub_255_2_n_1);
 assign sub_255_2_n_26 = ~(sub_255_2_n_18 | sub_255_2_n_17);
 assign sub_255_2_n_25 = ~(sub_255_2_n_8 | sub_255_2_n_6);
 assign sub_255_2_n_24 = ~(sub_255_2_n_5 | sub_255_2_n_4);
 assign sub_255_2_n_23 = ~(sub_255_2_n_16 & sub_255_2_n_19);
 assign sub_255_2_n_22 = ~(sub_255_2_n_14 & sub_255_2_n_20);
 assign sub_255_2_n_21 = ~(sub_255_2_n_7 | sub_255_2_n_9);
 assign sub_255_2_n_20 = ~({in2[10]} | {in2[11]});
 assign sub_255_2_n_19 = ~({in2[22]} | {in2[23]});
 assign sub_255_2_n_18 = ~(sub_255_2_n_11 | ~sub_255_2_n_13);
 assign sub_255_2_n_16 = ~({in2[20]} | {in2[21]});
 assign sub_255_2_n_15 = ~({in2[2]} | {in2[3]});
 assign sub_255_2_n_14 = ~({in2[8]} | {in2[9]});
 assign sub_255_2_n_17 = ~(in1_5_1_ | sub_255_2_n_13);
 assign sub_255_2_n_13 = ~{in2[2]};
 assign sub_255_2_n_12 = ~{in2[1]};
 assign sub_255_2_n_11 = ~in1_5_1_;
 assign sub_255_2_n_9 = ({in2[14]} | {in2[15]});
 assign sub_255_2_n_8 = ({in2[4]} | {in2[5]});
 assign sub_255_2_n_7 = ({in2[12]} | {in2[13]});
 assign sub_255_2_n_6 = ({in2[6]} | {in2[7]});
 assign sub_255_2_n_5 = ({in2[16]} | {in2[17]});
 assign sub_255_2_n_4 = ({in2[18]} | {in2[19]});
 assign sub_255_2_n_3 = (sub_255_2_n_1 & (in1_5_0_ | sub_255_2_n_12));
 assign sub_255_2_n_2 = ~({in1[46]} & ~{in2[0]});
 assign sub_255_2_n_1 = ~({in2[0]} & ~{in1[46]});
 assign sub_255_2_n_0 = (in1_5_0_ & sub_255_2_n_12);
 assign in1_10_24_ = ~(sub_274_2_n_42 & ~sub_274_2_n_33);
 assign in1_10_3_ = ~((sub_274_2_n_28 & ~sub_274_2_n_41) | (sub_274_2_n_29 & sub_274_2_n_41));
 assign sub_274_2_n_42 = ~(sub_274_2_n_30 & (sub_274_2_n_37 | sub_274_2_n_19));
 assign sub_274_2_n_41 = ~(sub_274_2_n_0 | ~(sub_274_2_n_36 | sub_274_2_n_14));
 assign in1_10_2_ = ~(sub_274_2_n_38 & ~sub_274_2_n_39);
 assign sub_274_2_n_39 = ~(sub_274_2_n_36 | sub_274_2_n_27);
 assign sub_274_2_n_38 = ~(sub_274_2_n_36 & sub_274_2_n_27);
 assign sub_274_2_n_37 = ~(sub_274_2_n_35 & ~sub_274_2_n_14);
 assign sub_274_2_n_36 = ~sub_274_2_n_35;
 assign sub_274_2_n_35 = ((sub_274_2_n_2 & in1_8_0_) | ((in1_8_0_ & sub_274_2_n_5) | (sub_274_2_n_5 &
    sub_274_2_n_2)));
 assign in1_10_1_ = (in1_8_0_ ^ (sub_274_2_n_5 ^ sub_274_2_n_2));
 assign sub_274_2_n_33 = ~(sub_274_2_n_32 & (sub_274_2_n_31 & ~sub_274_2_n_23));
 assign sub_274_2_n_32 = ~(sub_274_2_n_20 | sub_274_2_n_22);
 assign sub_274_2_n_31 = ~(sub_274_2_n_24 | sub_274_2_n_21);
 assign sub_274_2_n_30 = ~(sub_274_2_n_26 | sub_274_2_n_1);
 assign sub_274_2_n_29 = ~sub_274_2_n_28;
 assign sub_274_2_n_28 = ~(sub_274_2_n_1 | sub_274_2_n_19);
 assign sub_274_2_n_27 = ~(sub_274_2_n_0 | sub_274_2_n_14);
 assign sub_274_2_n_26 = ~(sub_274_2_n_19 | ~sub_274_2_n_0);
 assign in1_10_0_ = ~(sub_274_2_n_17 & sub_274_2_n_2);
 assign sub_274_2_n_24 = ~(sub_274_2_n_10 & sub_274_2_n_16);
 assign sub_274_2_n_23 = ~(sub_274_2_n_15 & sub_274_2_n_18);
 assign sub_274_2_n_22 = ~(sub_274_2_n_12 & sub_274_2_n_7);
 assign sub_274_2_n_21 = ~(sub_274_2_n_8 & sub_274_2_n_11);
 assign sub_274_2_n_20 = ~(sub_274_2_n_13 & sub_274_2_n_9);
 assign sub_274_2_n_18 = ~({in2[22]} | {in2[23]});
 assign sub_274_2_n_17 = ~({in1[45]} & ~{in2[0]});
 assign sub_274_2_n_16 = ~({in2[6]} | {in2[7]});
 assign sub_274_2_n_15 = ~({in2[20]} | {in2[21]});
 assign sub_274_2_n_19 = ~(in1_8_2_ | sub_274_2_n_4);
 assign sub_274_2_n_13 = ~({in2[8]} | {in2[9]});
 assign sub_274_2_n_12 = ~({in2[12]} | {in2[13]});
 assign sub_274_2_n_11 = ~({in2[18]} | {in2[19]});
 assign sub_274_2_n_10 = ~({in2[4]} | {in2[5]});
 assign sub_274_2_n_9 = ~({in2[10]} | {in2[11]});
 assign sub_274_2_n_8 = ~({in2[16]} | {in2[17]});
 assign sub_274_2_n_7 = ~({in2[14]} | {in2[15]});
 assign sub_274_2_n_14 = ~(in1_8_1_ | sub_274_2_n_6);
 assign sub_274_2_n_6 = ~{in2[2]};
 assign sub_274_2_n_5 = ~{in2[1]};
 assign sub_274_2_n_4 = ~{in2[3]};
 assign sub_274_2_n_2 = ~({in2[0]} & ~{in1[45]});
 assign sub_274_2_n_1 = (in1_8_2_ & sub_274_2_n_4);
 assign sub_274_2_n_0 = (in1_8_1_ & sub_274_2_n_6);
 assign in1_13_24_ = ~(sub_293_2_n_48 & (sub_293_2_n_49 | sub_293_2_n_30));
 assign in1_13_2_ = ~(sub_293_2_n_46 & ~sub_293_2_n_47);
 assign sub_293_2_n_50 = ~(sub_293_2_n_6 & ~(sub_293_2_n_44 & sub_293_2_n_38));
 assign sub_293_2_n_49 = ~(sub_293_2_n_42 & sub_293_2_n_12);
 assign sub_293_2_n_48 = ~(sub_293_2_n_43 | ~(sub_293_2_n_37 | sub_293_2_n_28));
 assign sub_293_2_n_47 = ~(sub_293_2_n_45 | sub_293_2_n_9);
 assign sub_293_2_n_46 = ~(sub_293_2_n_45 & sub_293_2_n_9);
 assign sub_293_2_n_45 = ~sub_293_2_n_44;
 assign sub_293_2_n_44 = ~((sub_293_2_n_0 & sub_293_2_n_14) | ((sub_293_2_n_14 & {in2[1]}) | ({in2[1]}
    & sub_293_2_n_0)));
 assign sub_293_2_n_43 = ~(sub_293_2_n_41 & sub_293_2_n_39);
 assign sub_293_2_n_42 = ~(sub_293_2_n_40 & sub_293_2_n_36);
 assign sub_293_2_n_41 = ~(sub_293_2_n_35 | (sub_293_2_n_34 | sub_293_2_n_31));
 assign sub_293_2_n_40 = ~(sub_293_2_n_0 & ~(sub_293_2_n_16 & in1_11_0_));
 assign sub_293_2_n_39 = ~(sub_293_2_n_32 | sub_293_2_n_33);
 assign sub_293_2_n_38 = ~(sub_293_2_n_4 | sub_293_2_n_3);
 assign sub_293_2_n_37 = ~(sub_293_2_n_3 | sub_293_2_n_23);
 assign sub_293_2_n_36 = ~(sub_293_2_n_4 | (sub_293_2_n_14 & {in2[1]}));
 assign sub_293_2_n_35 = ~(sub_293_2_n_25 & sub_293_2_n_18);
 assign sub_293_2_n_34 = ~(sub_293_2_n_20 & ~{in2[15]});
 assign sub_293_2_n_33 = ~(sub_293_2_n_27 & sub_293_2_n_26);
 assign sub_293_2_n_32 = ~(sub_293_2_n_17 & sub_293_2_n_24);
 assign sub_293_2_n_31 = ~(sub_293_2_n_21 & sub_293_2_n_19);
 assign sub_293_2_n_30 = ~(sub_293_2_n_22 & sub_293_2_n_29);
 assign sub_293_2_n_29 = ~sub_293_2_n_28;
 assign sub_293_2_n_27 = ~({in2[19]} | {in2[20]});
 assign sub_293_2_n_26 = ~({in2[21]} | {in2[22]});
 assign sub_293_2_n_25 = ~({in2[5]} | {in2[16]});
 assign sub_293_2_n_24 = ~({in2[9]} | {in2[10]});
 assign sub_293_2_n_28 = (sub_293_2_n_15 & in1_11_3_);
 assign sub_293_2_n_12 = ~(in1_11_1_ & ~{in2[2]});
 assign sub_293_2_n_21 = ~({in2[11]} | {in2[12]});
 assign sub_293_2_n_20 = ~({in2[6]} | {in2[7]});
 assign sub_293_2_n_19 = ~({in2[13]} | {in2[14]});
 assign sub_293_2_n_18 = ~({in2[17]} | {in2[18]});
 assign sub_293_2_n_17 = ~({in2[8]} | {in2[23]});
 assign sub_293_2_n_23 = ~(in1_11_3_ | sub_293_2_n_15);
 assign sub_293_2_n_22 = ~(in1_11_2_ & ~{in2[3]});
 assign sub_293_2_n_16 = ~{in2[1]};
 assign sub_293_2_n_15 = ~{in2[4]};
 assign sub_293_2_n_14 = ~in1_11_0_;
 assign in1_13_3_ = ~(sub_293_2_n_49 ^ sub_293_2_n_5);
 assign in1_13_4_ = ~(sub_293_2_n_50 ^ sub_293_2_n_7);
 assign sub_293_2_n_9 = ~(sub_293_2_n_4 | ~sub_293_2_n_12);
 assign in1_13_0_ = ~(sub_293_2_n_1 & ~sub_293_2_n_0);
 assign sub_293_2_n_7 = ~(sub_293_2_n_29 & ~sub_293_2_n_23);
 assign sub_293_2_n_6 = (sub_293_2_n_22 & (sub_293_2_n_12 | sub_293_2_n_3));
 assign sub_293_2_n_5 = ~(sub_293_2_n_22 & ~sub_293_2_n_3);
 assign sub_293_2_n_4 = ~(in1_11_1_ | ~{in2[2]});
 assign sub_293_2_n_3 = ~(in1_11_2_ | ~{in2[3]});
 assign in1_13_1_ = ~(sub_293_2_n_14 ^ ({in2[1]} ^ sub_293_2_n_0));
 assign sub_293_2_n_1 = ~({in1[44]} & ~{in2[0]});
 assign sub_293_2_n_0 = ~({in1[44]} | ~{in2[0]});
 assign in1_16_24_ = ~(sub_312_2_n_54 & sub_312_2_n_46);
 assign in1_16_5_ = ~(sub_312_2_n_55 & ~sub_312_2_n_56);
 assign in1_16_4_ = (sub_312_2_n_53 ^ sub_312_2_n_6);
 assign sub_312_2_n_56 = ~(sub_312_2_n_50 | sub_312_2_n_5);
 assign sub_312_2_n_55 = ~(sub_312_2_n_50 & sub_312_2_n_5);
 assign sub_312_2_n_54 = ~(sub_312_2_n_49 | sub_312_2_n_9);
 assign sub_312_2_n_53 = ~(sub_312_2_n_37 & ~(sub_312_2_n_47 & sub_312_2_n_33));
 assign sub_312_2_n_52 = ~(sub_312_2_n_26 | ~(sub_312_2_n_44 | sub_312_2_n_2));
 assign in1_16_2_ = ~((sub_312_2_n_44 & ~sub_312_2_n_34) | (sub_312_2_n_47 & sub_312_2_n_34));
 assign sub_312_2_n_50 = ~(sub_312_2_n_42 | (sub_312_2_n_48 | ~sub_312_2_n_24));
 assign sub_312_2_n_49 = ~(sub_312_2_n_43 | sub_312_2_n_7);
 assign sub_312_2_n_48 = ~(sub_312_2_n_39 | sub_312_2_n_44);
 assign sub_312_2_n_47 = ~sub_312_2_n_44;
 assign sub_312_2_n_46 = ~(sub_312_2_n_27 | (sub_312_2_n_45 | ~sub_312_2_n_29));
 assign sub_312_2_n_45 = ~(sub_312_2_n_40 & sub_312_2_n_28);
 assign sub_312_2_n_44 = ~(sub_312_2_n_41 | sub_312_2_n_14);
 assign sub_312_2_n_43 = ~(sub_312_2_n_37 & sub_312_2_n_38);
 assign sub_312_2_n_42 = ~(sub_312_2_n_37 | sub_312_2_n_3);
 assign sub_312_2_n_41 = ~(sub_312_2_n_15 | ~sub_312_2_n_23);
 assign sub_312_2_n_40 = ~(sub_312_2_n_31 | (sub_312_2_n_32 | ({in2[6]} | {in2[7]})));
 assign sub_312_2_n_39 = ~(sub_312_2_n_33 & ~sub_312_2_n_3);
 assign sub_312_2_n_38 = ~(sub_312_2_n_4 & ~(sub_312_2_n_24 & sub_312_2_n_19));
 assign sub_312_2_n_37 = ~(sub_312_2_n_35 | sub_312_2_n_1);
 assign sub_312_2_n_35 = ~(sub_312_2_n_25 | sub_312_2_n_18);
 assign sub_312_2_n_36 = ~(sub_312_2_n_1 | sub_312_2_n_18);
 assign sub_312_2_n_34 = ~(sub_312_2_n_26 | sub_312_2_n_2);
 assign sub_312_2_n_32 = ~(sub_312_2_n_16 & sub_312_2_n_17);
 assign sub_312_2_n_31 = ~(sub_312_2_n_20 & sub_312_2_n_21);
 assign in1_16_0_ = ~(sub_312_2_n_22 & sub_312_2_n_23);
 assign sub_312_2_n_29 = ~({in2[20]} | ({in2[21]} | ({in2[22]} | {in2[23]})));
 assign sub_312_2_n_28 = ~({in2[8]} | ({in2[9]} | ({in2[10]} | {in2[11]})));
 assign sub_312_2_n_33 = ~(sub_312_2_n_2 | sub_312_2_n_18);
 assign sub_312_2_n_27 = ~sub_312_2_n_4;
 assign sub_312_2_n_26 = ~sub_312_2_n_25;
 assign sub_312_2_n_22 = ~({in1[43]} & ~{in2[0]});
 assign sub_312_2_n_21 = ~({in2[14]} | {in2[15]});
 assign sub_312_2_n_20 = ~({in2[12]} | {in2[13]});
 assign sub_312_2_n_25 = ~(in1_14_1_ & ~{in2[2]});
 assign sub_312_2_n_24 = ~(in1_14_3_ & ~{in2[4]});
 assign sub_312_2_n_23 = ~({in2[0]} & ~{in1[43]});
 assign sub_312_2_n_17 = ~({in2[18]} | {in2[19]});
 assign sub_312_2_n_16 = ~({in2[16]} | {in2[17]});
 assign sub_312_2_n_15 = ~(in1_14_0_ | sub_312_2_n_12);
 assign sub_312_2_n_14 = ~(sub_312_2_n_11 | ~sub_312_2_n_12);
 assign sub_312_2_n_19 = ~(in1_14_4_ & ~{in2[5]});
 assign sub_312_2_n_18 = ~(in1_14_2_ | sub_312_2_n_13);
 assign sub_312_2_n_13 = ~{in2[3]};
 assign sub_312_2_n_12 = ~{in2[1]};
 assign sub_312_2_n_11 = ~in1_14_0_;
 assign sub_312_2_n_9 = (sub_312_2_n_3 & sub_312_2_n_19);
 assign in1_16_3_ = ~(sub_312_2_n_52 ^ sub_312_2_n_36);
 assign sub_312_2_n_7 = ~(sub_312_2_n_44 | ~sub_312_2_n_33);
 assign sub_312_2_n_6 = ~(sub_312_2_n_3 | ~sub_312_2_n_24);
 assign sub_312_2_n_5 = ~(sub_312_2_n_27 | ~sub_312_2_n_19);
 assign sub_312_2_n_4 = ~({in2[5]} & ~in1_14_4_);
 assign sub_312_2_n_3 = ~(in1_14_3_ | ~{in2[4]});
 assign sub_312_2_n_2 = ~(in1_14_1_ | ~{in2[2]});
 assign sub_312_2_n_1 = (in1_14_2_ & sub_312_2_n_13);
 assign in1_16_1_ = (sub_312_2_n_11 ^ ({in2[1]} ^ sub_312_2_n_23));
 assign in1_19_6_ = ~((sub_331_2_n_8 & ~sub_331_2_n_58) | (sub_331_2_n_36 & sub_331_2_n_58));
 assign in1_19_5_ = ~((sub_331_2_n_7 & ~sub_331_2_n_56) | (sub_331_2_n_30 & sub_331_2_n_56));
 assign sub_331_2_n_58 = ~(sub_331_2_n_53 | sub_331_2_n_40);
 assign in1_19_24_ = ~(sub_331_2_n_48 & (sub_331_2_n_51 | sub_331_2_n_45));
 assign sub_331_2_n_56 = ~(sub_331_2_n_10 & (sub_331_2_n_52 | sub_331_2_n_2));
 assign in1_19_4_ = ~((sub_331_2_n_6 & ~sub_331_2_n_52) | (sub_331_2_n_29 & sub_331_2_n_52));
 assign in1_19_3_ = ~(sub_331_2_n_50 ^ sub_331_2_n_32);
 assign sub_331_2_n_53 = ~(sub_331_2_n_38 | (sub_331_2_n_50 & sub_331_2_n_23));
 assign sub_331_2_n_52 = ~sub_331_2_n_51;
 assign sub_331_2_n_51 = ~(sub_331_2_n_9 & sub_331_2_n_39);
 assign sub_331_2_n_50 = ~(sub_331_2_n_49 | sub_331_2_n_16);
 assign sub_331_2_n_49 = ~(sub_331_2_n_46 | sub_331_2_n_3);
 assign sub_331_2_n_48 = ~(sub_331_2_n_47 | (sub_331_2_n_44 & sub_331_2_n_35));
 assign sub_331_2_n_47 = ~(sub_331_2_n_42 & (sub_331_2_n_37 | sub_331_2_n_33));
 assign sub_331_2_n_46 = ~(sub_331_2_n_43 | sub_331_2_n_20);
 assign sub_331_2_n_45 = ~sub_331_2_n_44;
 assign sub_331_2_n_44 = ~(sub_331_2_n_40 | sub_331_2_n_37);
 assign sub_331_2_n_43 = ~(sub_331_2_n_41 | ~(in1_17_0_ | sub_331_2_n_14));
 assign sub_331_2_n_42 = (sub_331_2_n_24 & (sub_331_2_n_25 & (sub_331_2_n_28 & sub_331_2_n_27)));
 assign sub_331_2_n_41 = ~sub_331_2_n_21;
 assign sub_331_2_n_40 = ~(sub_331_2_n_17 | (sub_331_2_n_10 & sub_331_2_n_18));
 assign sub_331_2_n_39 = ~(sub_331_2_n_22 | ~(sub_331_2_n_15 | sub_331_2_n_1));
 assign sub_331_2_n_38 = ~(sub_331_2_n_34 & ~(sub_331_2_n_1 & sub_331_2_n_23));
 assign sub_331_2_n_36 = ~sub_331_2_n_8;
 assign sub_331_2_n_35 = ~sub_331_2_n_34;
 assign sub_331_2_n_33 = ~(sub_331_2_n_5 | {in2[7]});
 assign sub_331_2_n_37 = ~(sub_331_2_n_19 | {in2[7]});
 assign sub_331_2_n_32 = ~(sub_331_2_n_22 | sub_331_2_n_1);
 assign sub_331_2_n_34 = ~(sub_331_2_n_2 | sub_331_2_n_17);
 assign sub_331_2_n_31 = ~(sub_331_2_n_16 | sub_331_2_n_3);
 assign sub_331_2_n_30 = ~sub_331_2_n_7;
 assign sub_331_2_n_29 = ~sub_331_2_n_6;
 assign sub_331_2_n_28 = ~({in2[16]} | ({in2[17]} | ({in2[18]} | {in2[19]})));
 assign sub_331_2_n_27 = ~({in2[20]} | ({in2[21]} | ({in2[22]} | {in2[23]})));
 assign in1_19_0_ = ~(sub_331_2_n_21 & ~(sub_331_2_n_12 & {in1[42]}));
 assign sub_331_2_n_25 = ~({in2[12]} | ({in2[13]} | ({in2[14]} | {in2[15]})));
 assign sub_331_2_n_24 = ~({in2[8]} | ({in2[9]} | ({in2[10]} | {in2[11]})));
 assign sub_331_2_n_22 = ~sub_331_2_n_23;
 assign sub_331_2_n_20 = ~(sub_331_2_n_13 | ~sub_331_2_n_14);
 assign sub_331_2_n_23 = ~(in1_17_2_ & ~{in2[3]});
 assign sub_331_2_n_21 = ~({in2[0]} & ~{in1[42]});
 assign sub_331_2_n_16 = ~sub_331_2_n_15;
 assign sub_331_2_n_19 = ~(in1_17_5_ & ~{in2[6]});
 assign sub_331_2_n_18 = ~(in1_17_4_ & ~{in2[5]});
 assign sub_331_2_n_17 = ~(in1_17_4_ | ~{in2[5]});
 assign sub_331_2_n_15 = ~(in1_17_1_ & ~{in2[2]});
 assign sub_331_2_n_10 = ~(in1_17_3_ & ~{in2[4]});
 assign sub_331_2_n_14 = ~{in2[1]};
 assign sub_331_2_n_13 = ~in1_17_0_;
 assign sub_331_2_n_12 = ~{in2[0]};
 assign sub_331_2_n_9 = ~(sub_331_2_n_49 & ~sub_331_2_n_1);
 assign sub_331_2_n_8 = ~(sub_331_2_n_5 | ~sub_331_2_n_19);
 assign sub_331_2_n_7 = ~(sub_331_2_n_18 & ~sub_331_2_n_17);
 assign sub_331_2_n_6 = ~(sub_331_2_n_2 | ~sub_331_2_n_10);
 assign sub_331_2_n_5 = ~(in1_17_5_ | ~{in2[6]});
 assign sub_331_2_n_3 = ~(in1_17_1_ | ~{in2[2]});
 assign sub_331_2_n_2 = ~(in1_17_3_ | ~{in2[4]});
 assign sub_331_2_n_1 = ~(in1_17_2_ | ~{in2[3]});
 assign in1_19_2_ = ~(sub_331_2_n_31 ^ sub_331_2_n_46);
 assign in1_19_1_ = (sub_331_2_n_13 ^ ({in2[1]} ^ sub_331_2_n_21));
 assign in1_22_6_ = ~((sub_350_2_n_50 & ~sub_350_2_n_78) | (sub_350_2_n_49 & sub_350_2_n_78));
 assign sub_350_2_n_82 = ~(sub_350_2_n_14 & (sub_350_2_n_74 | sub_350_2_n_9));
 assign in1_22_24_ = ~(sub_350_2_n_68 & (sub_350_2_n_73 | sub_350_2_n_61));
 assign in1_22_4_ = ~((sub_350_2_n_7 & ~sub_350_2_n_75) | (sub_350_2_n_43 & sub_350_2_n_75));
 assign sub_350_2_n_79 = ~(sub_350_2_n_66 & (sub_350_2_n_75 | sub_350_2_n_57));
 assign sub_350_2_n_78 = ~(sub_350_2_n_65 & sub_350_2_n_76);
 assign in1_22_3_ = ~((sub_350_2_n_5 & ~sub_350_2_n_71) | (sub_350_2_n_40 & sub_350_2_n_71));
 assign sub_350_2_n_76 = ~(sub_350_2_n_69 & sub_350_2_n_39);
 assign sub_350_2_n_75 = ~(sub_350_2_n_69 | sub_350_2_n_56);
 assign sub_350_2_n_74 = ~(sub_350_2_n_70 | sub_350_2_n_48);
 assign sub_350_2_n_73 = ~(sub_350_2_n_72 | sub_350_2_n_53);
 assign sub_350_2_n_72 = ~(sub_350_2_n_63 | sub_350_2_n_48);
 assign sub_350_2_n_71 = ~(sub_350_2_n_63 | sub_350_2_n_16);
 assign sub_350_2_n_70 = ~(sub_350_2_n_67 | sub_350_2_n_0);
 assign sub_350_2_n_69 = ~(sub_350_2_n_67 | sub_350_2_n_6);
 assign sub_350_2_n_68 = ~(sub_350_2_n_59 | (sub_350_2_n_52 & sub_350_2_n_8));
 assign sub_350_2_n_67 = ~(sub_350_2_n_60 | sub_350_2_n_4);
 assign sub_350_2_n_66 = ~(sub_350_2_n_26 | ~(sub_350_2_n_51 | sub_350_2_n_30));
 assign sub_350_2_n_65 = ~(sub_350_2_n_58 | ~sub_350_2_n_51);
 assign in1_22_1_ = ~(in1_20_0_ ^ ({in2[1]} ^ sub_350_2_n_28));
 assign sub_350_2_n_63 = ~(sub_350_2_n_62 | sub_350_2_n_10);
 assign sub_350_2_n_62 = ~(sub_350_2_n_28 | (sub_350_2_n_20 & in1_20_0_));
 assign sub_350_2_n_61 = ~(sub_350_2_n_51 & sub_350_2_n_52);
 assign sub_350_2_n_60 = ~(sub_350_2_n_23 | ~sub_350_2_n_28);
 assign sub_350_2_n_59 = ~(sub_350_2_n_35 & (sub_350_2_n_36 & (sub_350_2_n_34 & sub_350_2_n_38)));
 assign sub_350_2_n_58 = ~(sub_350_2_n_54 & sub_350_2_n_55);
 assign sub_350_2_n_57 = ~(sub_350_2_n_39 & ~sub_350_2_n_30);
 assign sub_350_2_n_56 = ~(sub_350_2_n_24 & (sub_350_2_n_31 | sub_350_2_n_3));
 assign sub_350_2_n_55 = ~(sub_350_2_n_39 & ~sub_350_2_n_24);
 assign sub_350_2_n_54 = ~(sub_350_2_n_44 & sub_350_2_n_39);
 assign sub_350_2_n_53 = ~(sub_350_2_n_41 & sub_350_2_n_39);
 assign sub_350_2_n_52 = ~(sub_350_2_n_45 | sub_350_2_n_1);
 assign sub_350_2_n_51 = ~(sub_350_2_n_33 | ~(sub_350_2_n_14 | sub_350_2_n_32));
 assign sub_350_2_n_50 = ~sub_350_2_n_49;
 assign sub_350_2_n_45 = ~(sub_350_2_n_25 | sub_350_2_n_15);
 assign sub_350_2_n_44 = ~(sub_350_2_n_3 | ~sub_350_2_n_16);
 assign sub_350_2_n_49 = ~(sub_350_2_n_26 | sub_350_2_n_30);
 assign sub_350_2_n_48 = ~(sub_350_2_n_31 & sub_350_2_n_24);
 assign sub_350_2_n_47 = ~(sub_350_2_n_16 | sub_350_2_n_0);
 assign sub_350_2_n_46 = ~(sub_350_2_n_1 | sub_350_2_n_15);
 assign sub_350_2_n_43 = ~sub_350_2_n_7;
 assign sub_350_2_n_40 = ~sub_350_2_n_5;
 assign sub_350_2_n_38 = ~({in2[20]} | ({in2[21]} | ({in2[22]} | {in2[23]})));
 assign in1_22_0_ = ~(sub_350_2_n_28 & ~(sub_350_2_n_21 & {in1[41]}));
 assign sub_350_2_n_36 = ~({in2[12]} | ({in2[13]} | ({in2[14]} | {in2[15]})));
 assign sub_350_2_n_35 = ~({in2[8]} | ({in2[9]} | ({in2[10]} | {in2[11]})));
 assign sub_350_2_n_34 = ~({in2[16]} | ({in2[17]} | ({in2[18]} | {in2[19]})));
 assign sub_350_2_n_42 = ~(sub_350_2_n_33 | sub_350_2_n_32);
 assign sub_350_2_n_41 = ~(sub_350_2_n_3 & sub_350_2_n_24);
 assign sub_350_2_n_39 = ~(sub_350_2_n_2 | sub_350_2_n_32);
 assign sub_350_2_n_31 = ~sub_350_2_n_16;
 assign sub_350_2_n_30 = ~sub_350_2_n_29;
 assign sub_350_2_n_27 = (in1_20_0_ | sub_350_2_n_20);
 assign sub_350_2_n_33 = (sub_350_2_n_22 & in1_20_4_);
 assign sub_350_2_n_32 = ~(in1_20_4_ | sub_350_2_n_22);
 assign sub_350_2_n_16 = ~({in2[2]} | ~in1_20_1_);
 assign sub_350_2_n_29 = ~(sub_350_2_n_18 & {in2[6]});
 assign sub_350_2_n_28 = ~({in2[0]} & ~{in1[41]});
 assign sub_350_2_n_26 = ~sub_350_2_n_25;
 assign sub_350_2_n_23 = ~(in1_20_0_ | sub_350_2_n_20);
 assign sub_350_2_n_25 = ~(in1_20_5_ & ~{in2[6]});
 assign sub_350_2_n_15 = ~(in1_20_6_ | sub_350_2_n_19);
 assign sub_350_2_n_14 = ~(in1_20_3_ & ~{in2[4]});
 assign sub_350_2_n_24 = ~(in1_20_2_ & ~{in2[3]});
 assign sub_350_2_n_22 = ~{in2[5]};
 assign sub_350_2_n_21 = ~{in2[0]};
 assign sub_350_2_n_20 = ~{in2[1]};
 assign sub_350_2_n_19 = ~{in2[7]};
 assign sub_350_2_n_18 = ~in1_20_5_;
 assign in1_22_2_ = ~(sub_350_2_n_67 ^ sub_350_2_n_47);
 assign in1_22_7_ = (sub_350_2_n_79 ^ sub_350_2_n_46);
 assign in1_22_5_ = (sub_350_2_n_82 ^ sub_350_2_n_42);
 assign sub_350_2_n_10 = ~(sub_350_2_n_27 & ~sub_350_2_n_0);
 assign sub_350_2_n_9 = ~(sub_350_2_n_41 & ~sub_350_2_n_2);
 assign sub_350_2_n_8 = ~(sub_350_2_n_29 & ~sub_350_2_n_15);
 assign sub_350_2_n_7 = ~(sub_350_2_n_2 | ~sub_350_2_n_14);
 assign sub_350_2_n_6 = (sub_350_2_n_3 | sub_350_2_n_0);
 assign sub_350_2_n_5 = ~(sub_350_2_n_3 | ~sub_350_2_n_24);
 assign sub_350_2_n_4 = (in1_20_0_ & sub_350_2_n_20);
 assign sub_350_2_n_3 = ~(in1_20_2_ | ~{in2[3]});
 assign sub_350_2_n_2 = ~(in1_20_3_ | ~{in2[4]});
 assign sub_350_2_n_1 = (in1_20_6_ & sub_350_2_n_19);
 assign sub_350_2_n_0 = ~(in1_20_1_ | ~{in2[2]});
 assign in1_25_8_ = (sub_369_2_n_86 ^ sub_369_2_n_42);
 assign in1_25_7_ = (sub_369_2_n_85 ^ sub_369_2_n_7);
 assign in1_25_4_ = (sub_369_2_n_79 ^ sub_369_2_n_8);
 assign sub_369_2_n_86 = ~(sub_369_2_n_69 | (sub_369_2_n_79 & sub_369_2_n_58));
 assign sub_369_2_n_85 = ~(sub_369_2_n_67 & ~(sub_369_2_n_79 & sub_369_2_n_57));
 assign sub_369_2_n_84 = ~(sub_369_2_n_33 & (sub_369_2_n_13 | sub_369_2_n_6));
 assign in1_25_24_ = ~sub_369_2_n_82;
 assign sub_369_2_n_82 = ~(sub_369_2_n_80 | sub_369_2_n_78);
 assign sub_369_2_n_81 = ~(sub_369_2_n_76 | sub_369_2_n_55);
 assign sub_369_2_n_80 = ~(sub_369_2_n_71 | sub_369_2_n_76);
 assign sub_369_2_n_79 = ~(sub_369_2_n_52 & (sub_369_2_n_72 | sub_369_2_n_0));
 assign sub_369_2_n_78 = ~(sub_369_2_n_59 & (sub_369_2_n_65 | sub_369_2_n_63));
 assign in1_25_2_ = ~(sub_369_2_n_74 & ~sub_369_2_n_73);
 assign sub_369_2_n_76 = ~(sub_369_2_n_75 | sub_369_2_n_51);
 assign sub_369_2_n_75 = ~(sub_369_2_n_64 | sub_369_2_n_50);
 assign sub_369_2_n_74 = ~(sub_369_2_n_68 & sub_369_2_n_41);
 assign sub_369_2_n_73 = ~(sub_369_2_n_68 | sub_369_2_n_41);
 assign sub_369_2_n_72 = ~(sub_369_2_n_68 & sub_369_2_n_1);
 assign sub_369_2_n_71 = ~(sub_369_2_n_70 & sub_369_2_n_56);
 assign sub_369_2_n_70 = ~(sub_369_2_n_63 | sub_369_2_n_55);
 assign sub_369_2_n_69 = ~(sub_369_2_n_56 & (sub_369_2_n_54 | sub_369_2_n_49));
 assign sub_369_2_n_68 = ~((sub_369_2_n_60 & sub_369_2_n_18) | ((sub_369_2_n_18 & {in2[1]}) | ({in2[1]}
    & sub_369_2_n_60)));
 assign sub_369_2_n_67 = ~(sub_369_2_n_26 | (sub_369_2_n_55 & sub_369_2_n_22));
 assign in1_25_1_ = ~(in1_23_0_ ^ (sub_369_2_n_19 ^ sub_369_2_n_60));
 assign sub_369_2_n_65 = ~(sub_369_2_n_44 | (sub_369_2_n_62 | ~sub_369_2_n_30));
 assign sub_369_2_n_64 = ~(sub_369_2_n_61 | sub_369_2_n_45);
 assign sub_369_2_n_63 = ~(sub_369_2_n_28 | ~sub_369_2_n_53);
 assign sub_369_2_n_62 = ~(sub_369_2_n_53 & (in1_23_7_ | sub_369_2_n_15));
 assign sub_369_2_n_61 = ~(sub_369_2_n_29 | (sub_369_2_n_19 & in1_23_0_));
 assign sub_369_2_n_60 = ~sub_369_2_n_29;
 assign sub_369_2_n_59 = (sub_369_2_n_36 & sub_369_2_n_37);
 assign sub_369_2_n_58 = ~(sub_369_2_n_47 | sub_369_2_n_49);
 assign sub_369_2_n_57 = ~(sub_369_2_n_47 | sub_369_2_n_2);
 assign sub_369_2_n_56 = ~(sub_369_2_n_43 & sub_369_2_n_30);
 assign sub_369_2_n_54 = ~sub_369_2_n_55;
 assign sub_369_2_n_55 = ~(sub_369_2_n_4 | (sub_369_2_n_33 & sub_369_2_n_34));
 assign sub_369_2_n_53 = ~({in2[10]} | ({in2[11]} | ({in2[15]} | sub_369_2_n_35)));
 assign sub_369_2_n_52 = ~(sub_369_2_n_32 | ~(sub_369_2_n_23 | sub_369_2_n_0));
 assign sub_369_2_n_51 = ~(sub_369_2_n_39 & sub_369_2_n_46);
 assign sub_369_2_n_47 = ~sub_369_2_n_46;
 assign sub_369_2_n_45 = ~(sub_369_2_n_1 & ~sub_369_2_n_21);
 assign sub_369_2_n_44 = ~(sub_369_2_n_3 | ~sub_369_2_n_2);
 assign sub_369_2_n_43 = ~(sub_369_2_n_25 & sub_369_2_n_27);
 assign sub_369_2_n_50 = ~(sub_369_2_n_23 & sub_369_2_n_31);
 assign sub_369_2_n_42 = ~(sub_369_2_n_28 & ~(sub_369_2_n_20 & {in2[8]}));
 assign sub_369_2_n_49 = ~(sub_369_2_n_30 & ~sub_369_2_n_2);
 assign sub_369_2_n_48 = ~(sub_369_2_n_32 | sub_369_2_n_0);
 assign sub_369_2_n_46 = ~(sub_369_2_n_24 | sub_369_2_n_4);
 assign sub_369_2_n_39 = ~(sub_369_2_n_0 & sub_369_2_n_31);
 assign in1_25_0_ = ~(sub_369_2_n_29 & ~(sub_369_2_n_17 & {in1[40]}));
 assign sub_369_2_n_37 = ~({in2[20]} | ({in2[21]} | ({in2[22]} | {in2[23]})));
 assign sub_369_2_n_36 = ~({in2[16]} | ({in2[17]} | ({in2[18]} | {in2[19]})));
 assign sub_369_2_n_35 = ({in2[9]} | ({in2[12]} | ({in2[13]} | {in2[14]})));
 assign sub_369_2_n_41 = ~(sub_369_2_n_23 & sub_369_2_n_1);
 assign sub_369_2_n_40 = ~(sub_369_2_n_26 | sub_369_2_n_2);
 assign sub_369_2_n_32 = ~sub_369_2_n_31;
 assign sub_369_2_n_34 = ~(in1_23_4_ & ~{in2[5]});
 assign sub_369_2_n_33 = ~(in1_23_3_ & ~{in2[4]});
 assign sub_369_2_n_31 = ~(in1_23_2_ & ~{in2[3]});
 assign sub_369_2_n_30 = ~(sub_369_2_n_16 & {in2[7]});
 assign sub_369_2_n_29 = ({in1[40]} | sub_369_2_n_17);
 assign sub_369_2_n_27 = ~sub_369_2_n_3;
 assign sub_369_2_n_26 = ~sub_369_2_n_25;
 assign sub_369_2_n_22 = ~sub_369_2_n_2;
 assign sub_369_2_n_28 = ~(in1_23_7_ & ~{in2[8]});
 assign sub_369_2_n_21 = ~(in1_23_0_ | sub_369_2_n_19);
 assign sub_369_2_n_25 = ~(in1_23_5_ & ~{in2[6]});
 assign sub_369_2_n_24 = ~(in1_23_3_ | ~{in2[4]});
 assign sub_369_2_n_23 = ~(in1_23_1_ & ~{in2[2]});
 assign sub_369_2_n_20 = ~in1_23_7_;
 assign sub_369_2_n_19 = ~{in2[1]};
 assign sub_369_2_n_18 = ~in1_23_0_;
 assign sub_369_2_n_17 = ~{in2[0]};
 assign sub_369_2_n_16 = ~in1_23_6_;
 assign sub_369_2_n_15 = ~{in2[8]};
 assign sub_369_2_n_13 = ~(sub_369_2_n_50 | ~sub_369_2_n_72);
 assign in1_25_3_ = ~(sub_369_2_n_5 ^ sub_369_2_n_48);
 assign in1_25_5_ = (sub_369_2_n_84 ^ sub_369_2_n_9);
 assign in1_25_6_ = ~(sub_369_2_n_81 ^ sub_369_2_n_40);
 assign sub_369_2_n_9 = ~(sub_369_2_n_4 | ~sub_369_2_n_34);
 assign sub_369_2_n_8 = ~(sub_369_2_n_24 | ~sub_369_2_n_33);
 assign sub_369_2_n_7 = ~(sub_369_2_n_3 | ~sub_369_2_n_30);
 assign sub_369_2_n_6 = (sub_369_2_n_0 | sub_369_2_n_24);
 assign sub_369_2_n_5 = ~(sub_369_2_n_64 | ~sub_369_2_n_23);
 assign sub_369_2_n_4 = ~(in1_23_4_ | ~{in2[5]});
 assign sub_369_2_n_3 = ~(sub_369_2_n_16 | {in2[7]});
 assign sub_369_2_n_2 = ~(in1_23_5_ | ~{in2[6]});
 assign sub_369_2_n_1 = ~({in2[2]} & ~in1_23_1_);
 assign sub_369_2_n_0 = ~(in1_23_2_ | ~{in2[3]});
 assign in1_28_9_ = ~(~(sub_388_2_n_110 & sub_388_2_n_10) & (sub_388_2_n_110 | sub_388_2_n_10));
 assign sub_388_2_n_110 = ~(sub_388_2_n_20 & (sub_388_2_n_107 | sub_388_2_n_7));
 assign in1_28_24_ = ~(sub_388_2_n_108 & sub_388_2_n_98);
 assign sub_388_2_n_108 = ~(sub_388_2_n_104 & sub_388_2_n_86);
 assign sub_388_2_n_107 = ~(sub_388_2_n_100 | sub_388_2_n_85);
 assign sub_388_2_n_106 = ~(sub_388_2_n_38 | (sub_388_2_n_94 & sub_388_2_n_41));
 assign in1_28_4_ = ~(sub_388_2_n_94 ^ sub_388_2_n_44);
 assign sub_388_2_n_104 = ~(sub_388_2_n_103 & sub_388_2_n_76);
 assign sub_388_2_n_103 = ~(sub_388_2_n_93 & sub_388_2_n_63);
 assign sub_388_2_n_102 = ~(sub_388_2_n_87 & sub_388_2_n_96);
 assign sub_388_2_n_101 = ~(sub_388_2_n_97 | sub_388_2_n_72);
 assign sub_388_2_n_100 = ~(sub_388_2_n_71 | sub_388_2_n_99);
 assign sub_388_2_n_99 = ~(sub_388_2_n_92 | sub_388_2_n_30);
 assign sub_388_2_n_98 = ~(sub_388_2_n_70 | (sub_388_2_n_80 & sub_388_2_n_84));
 assign sub_388_2_n_97 = ~(sub_388_2_n_91 | sub_388_2_n_68);
 assign sub_388_2_n_96 = ~(sub_388_2_n_92 & sub_388_2_n_75);
 assign in1_28_2_ = ~(sub_388_2_n_90 & ~sub_388_2_n_89);
 assign sub_388_2_n_94 = ~sub_388_2_n_93;
 assign sub_388_2_n_93 = ~(sub_388_2_n_88 | sub_388_2_n_62);
 assign sub_388_2_n_91 = ~sub_388_2_n_92;
 assign sub_388_2_n_92 = ~(sub_388_2_n_82 & sub_388_2_n_36);
 assign sub_388_2_n_90 = ~(sub_388_2_n_83 & sub_388_2_n_11);
 assign sub_388_2_n_89 = ~(sub_388_2_n_83 | sub_388_2_n_11);
 assign sub_388_2_n_88 = ~(sub_388_2_n_83 | sub_388_2_n_55);
 assign sub_388_2_n_87 = ~(sub_388_2_n_73 | (sub_388_2_n_74 | ~sub_388_2_n_42));
 assign sub_388_2_n_86 = ~(sub_388_2_n_81 | sub_388_2_n_77);
 assign sub_388_2_n_85 = ~(sub_388_2_n_63 & (sub_388_2_n_61 | sub_388_2_n_58));
 assign sub_388_2_n_84 = ~(sub_388_2_n_79 & sub_388_2_n_40);
 assign sub_388_2_n_83 = ~(sub_388_2_n_78 | sub_388_2_n_29);
 assign sub_388_2_n_82 = ~(sub_388_2_n_18 & sub_388_2_n_50);
 assign sub_388_2_n_81 = ~sub_388_2_n_80;
 assign sub_388_2_n_79 = ~(sub_388_2_n_7 | ~sub_388_2_n_65);
 assign sub_388_2_n_78 = ~(sub_388_2_n_33 | ~sub_388_2_n_31);
 assign sub_388_2_n_77 = ~(sub_388_2_n_61 | sub_388_2_n_58);
 assign sub_388_2_n_80 = ~(sub_388_2_n_65 & (sub_388_2_n_52 | sub_388_2_n_8));
 assign sub_388_2_n_76 = ~(sub_388_2_n_66 & sub_388_2_n_63);
 assign sub_388_2_n_75 = ~(sub_388_2_n_64 | sub_388_2_n_5);
 assign sub_388_2_n_74 = ~(sub_388_2_n_64 | sub_388_2_n_19);
 assign sub_388_2_n_73 = ~(sub_388_2_n_61 | ~sub_388_2_n_32);
 assign sub_388_2_n_72 = ~(sub_388_2_n_69 & sub_388_2_n_61);
 assign sub_388_2_n_71 = ~(sub_388_2_n_67 & sub_388_2_n_49);
 assign sub_388_2_n_70 = ~(sub_388_2_n_46 & sub_388_2_n_47);
 assign sub_388_2_n_69 = ~(sub_388_2_n_56 & sub_388_2_n_30);
 assign sub_388_2_n_68 = ~(sub_388_2_n_56 & sub_388_2_n_21);
 assign sub_388_2_n_67 = ~sub_388_2_n_66;
 assign sub_388_2_n_66 = ~(sub_388_2_n_56 & sub_388_2_n_57);
 assign sub_388_2_n_65 = ~({in2[14]} | ({in2[15]} | ~sub_388_2_n_48));
 assign sub_388_2_n_64 = ~(sub_388_2_n_56 & sub_388_2_n_32);
 assign sub_388_2_n_63 = ~(sub_388_2_n_53 | sub_388_2_n_1);
 assign sub_388_2_n_62 = ~(sub_388_2_n_19 & (sub_388_2_n_36 | sub_388_2_n_5));
 assign sub_388_2_n_61 = ~(sub_388_2_n_54 | sub_388_2_n_6);
 assign sub_388_2_n_58 = ~sub_388_2_n_57;
 assign sub_388_2_n_55 = ~(sub_388_2_n_34 & sub_388_2_n_21);
 assign sub_388_2_n_54 = ~(sub_388_2_n_37 | sub_388_2_n_35);
 assign sub_388_2_n_53 = ~(sub_388_2_n_42 | sub_388_2_n_43);
 assign sub_388_2_n_52 = ~(sub_388_2_n_20 | sub_388_2_n_39);
 assign sub_388_2_n_60 = ~(sub_388_2_n_30 | sub_388_2_n_5);
 assign sub_388_2_n_59 = ~(sub_388_2_n_6 | sub_388_2_n_35);
 assign sub_388_2_n_57 = ~(sub_388_2_n_2 | sub_388_2_n_43);
 assign sub_388_2_n_56 = ~(sub_388_2_n_4 | sub_388_2_n_35);
 assign sub_388_2_n_50 = ~(sub_388_2_n_33 | sub_388_2_n_0);
 assign sub_388_2_n_49 = ~(sub_388_2_n_5 & sub_388_2_n_19);
 assign sub_388_2_n_48 = ~({in2[10]} | ({in2[11]} | ({in2[12]} | {in2[13]})));
 assign sub_388_2_n_47 = ~({in2[20]} | ({in2[21]} | ({in2[22]} | {in2[23]})));
 assign sub_388_2_n_46 = ~({in2[16]} | ({in2[17]} | ({in2[18]} | {in2[19]})));
 assign in1_28_0_ = ~(sub_388_2_n_31 & ~(sub_388_2_n_27 & {in1[39]}));
 assign sub_388_2_n_51 = ~(sub_388_2_n_1 | sub_388_2_n_43);
 assign sub_388_2_n_44 = ~(sub_388_2_n_37 & sub_388_2_n_41);
 assign sub_388_2_n_41 = ~sub_388_2_n_4;
 assign sub_388_2_n_40 = ~sub_388_2_n_39;
 assign sub_388_2_n_38 = ~sub_388_2_n_37;
 assign sub_388_2_n_21 = ~sub_388_2_n_5;
 assign sub_388_2_n_43 = ~(in1_26_6_ | sub_388_2_n_24);
 assign sub_388_2_n_42 = ~(in1_26_5_ & ~{in2[6]});
 assign sub_388_2_n_39 = ~(in1_26_8_ | sub_388_2_n_26);
 assign sub_388_2_n_37 = ~(in1_26_3_ & ~{in2[4]});
 assign sub_388_2_n_36 = ~(in1_26_1_ & ~{in2[2]});
 assign sub_388_2_n_35 = ~(in1_26_4_ | sub_388_2_n_23);
 assign sub_388_2_n_34 = ~sub_388_2_n_0;
 assign sub_388_2_n_32 = ~sub_388_2_n_2;
 assign sub_388_2_n_30 = ~sub_388_2_n_19;
 assign sub_388_2_n_29 = ~(sub_388_2_n_28 | ~sub_388_2_n_25);
 assign sub_388_2_n_33 = ~(in1_26_0_ | sub_388_2_n_25);
 assign sub_388_2_n_20 = ~(in1_26_7_ & ~{in2[8]});
 assign sub_388_2_n_31 = ~({in2[0]} & ~{in1[39]});
 assign sub_388_2_n_19 = ~(in1_26_2_ & ~{in2[3]});
 assign sub_388_2_n_28 = ~in1_26_0_;
 assign sub_388_2_n_27 = ~{in2[0]};
 assign sub_388_2_n_26 = ~{in2[9]};
 assign sub_388_2_n_25 = ~{in2[1]};
 assign sub_388_2_n_24 = ~{in2[7]};
 assign sub_388_2_n_23 = ~{in2[5]};
 assign sub_388_2_n_18 = (sub_388_2_n_31 | (sub_388_2_n_25 & in1_26_0_));
 assign in1_28_3_ = ~(sub_388_2_n_91 ^ sub_388_2_n_60);
 assign in1_28_6_ = ~(sub_388_2_n_101 ^ sub_388_2_n_12);
 assign in1_28_5_ = ~(sub_388_2_n_106 ^ sub_388_2_n_59);
 assign in1_28_8_ = ~(sub_388_2_n_107 ^ sub_388_2_n_9);
 assign in1_28_7_ = (sub_388_2_n_102 ^ sub_388_2_n_51);
 assign sub_388_2_n_12 = ~(sub_388_2_n_2 | ~sub_388_2_n_42);
 assign sub_388_2_n_11 = ~(sub_388_2_n_0 | ~sub_388_2_n_36);
 assign sub_388_2_n_10 = ~(sub_388_2_n_40 & ~sub_388_2_n_8);
 assign sub_388_2_n_9 = ~(sub_388_2_n_7 | ~sub_388_2_n_20);
 assign sub_388_2_n_8 = (in1_26_8_ & sub_388_2_n_26);
 assign sub_388_2_n_7 = ~(in1_26_7_ | ~{in2[8]});
 assign sub_388_2_n_6 = (in1_26_4_ & sub_388_2_n_23);
 assign sub_388_2_n_5 = ~(in1_26_2_ | ~{in2[3]});
 assign sub_388_2_n_4 = ~(in1_26_3_ | ~{in2[4]});
 assign sub_388_2_n_2 = ~(in1_26_5_ | ~{in2[6]});
 assign sub_388_2_n_1 = (in1_26_6_ & sub_388_2_n_24);
 assign sub_388_2_n_0 = ~(in1_26_1_ | ~{in2[2]});
 assign in1_28_1_ = (sub_388_2_n_28 ^ ({in2[1]} ^ sub_388_2_n_31));
 assign in1_31_10_ = ~((sub_407_2_n_57 & ~sub_407_2_n_86) | (sub_407_2_n_16 & sub_407_2_n_86));
 assign in1_31_9_ = ~((sub_407_2_n_52 & ~sub_407_2_n_89) | (sub_407_2_n_51 & sub_407_2_n_89));
 assign sub_407_2_n_89 = ~(sub_407_2_n_36 & (sub_407_2_n_83 | sub_407_2_n_6));
 assign in1_31_24_ = ~(sub_407_2_n_85 & sub_407_2_n_76);
 assign in1_31_8_ = ~(sub_407_2_n_83 ^ sub_407_2_n_11);
 assign sub_407_2_n_86 = ~(sub_407_2_n_66 & (sub_407_2_n_83 | sub_407_2_n_56));
 assign sub_407_2_n_85 = ~(sub_407_2_n_83 & sub_407_2_n_71);
 assign sub_407_2_n_84 = ~(sub_407_2_n_25 & (sub_407_2_n_82 | sub_407_2_n_4));
 assign sub_407_2_n_83 = ~(sub_407_2_n_19 | sub_407_2_n_75);
 assign sub_407_2_n_82 = ~(sub_407_2_n_62 | (sub_407_2_n_79 & sub_407_2_n_61));
 assign sub_407_2_n_81 = ~(sub_407_2_n_43 | (sub_407_2_n_79 & sub_407_2_n_2));
 assign sub_407_2_n_80 = ~(sub_407_2_n_39 & (sub_407_2_n_74 | sub_407_2_n_38));
 assign sub_407_2_n_79 = ~sub_407_2_n_78;
 assign sub_407_2_n_78 = ~(sub_407_2_n_77 | sub_407_2_n_64);
 assign sub_407_2_n_77 = ~(sub_407_2_n_53 | sub_407_2_n_74);
 assign sub_407_2_n_76 = ~(sub_407_2_n_69 | sub_407_2_n_65);
 assign sub_407_2_n_75 = ~(sub_407_2_n_72 & sub_407_2_n_63);
 assign sub_407_2_n_74 = ~(sub_407_2_n_70 | sub_407_2_n_0);
 assign in1_31_1_ = ~(in1_29_0_ ^ ({in2[1]} ^ sub_407_2_n_34));
 assign sub_407_2_n_72 = ~(sub_407_2_n_62 & sub_407_2_n_50);
 assign sub_407_2_n_71 = ~(sub_407_2_n_59 & (sub_407_2_n_58 | sub_407_2_n_60));
 assign sub_407_2_n_70 = ~(sub_407_2_n_33 | ~sub_407_2_n_34);
 assign sub_407_2_n_69 = ~(sub_407_2_n_68 & ~sub_407_2_n_67);
 assign sub_407_2_n_68 = ~(sub_407_2_n_5 | ~sub_407_2_n_47);
 assign sub_407_2_n_67 = ~(sub_407_2_n_45 & sub_407_2_n_48);
 assign sub_407_2_n_66 = ~(sub_407_2_n_58 | sub_407_2_n_41);
 assign sub_407_2_n_65 = ~(sub_407_2_n_60 | sub_407_2_n_55);
 assign sub_407_2_n_64 = ~(sub_407_2_n_54 & sub_407_2_n_7);
 assign sub_407_2_n_63 = ~(sub_407_2_n_9 | ~(sub_407_2_n_25 | sub_407_2_n_35));
 assign sub_407_2_n_62 = ~(sub_407_2_n_44 & (sub_407_2_n_42 | sub_407_2_n_3));
 assign sub_407_2_n_61 = ~sub_407_2_n_10;
 assign sub_407_2_n_59 = ~sub_407_2_n_5;
 assign sub_407_2_n_57 = ~sub_407_2_n_16;
 assign sub_407_2_n_56 = ~sub_407_2_n_55;
 assign sub_407_2_n_54 = ~(sub_407_2_n_40 & ~sub_407_2_n_39);
 assign sub_407_2_n_53 = ~(sub_407_2_n_40 & ~sub_407_2_n_38);
 assign sub_407_2_n_60 = ~(sub_407_2_n_37 & ~sub_407_2_n_41);
 assign sub_407_2_n_58 = ~(sub_407_2_n_36 | sub_407_2_n_1);
 assign sub_407_2_n_55 = ~(sub_407_2_n_6 | sub_407_2_n_1);
 assign sub_407_2_n_52 = ~sub_407_2_n_51;
 assign sub_407_2_n_48 = ~({in2[16]} | ({in2[17]} | ({in2[18]} | {in2[19]})));
 assign sub_407_2_n_47 = ~({in2[20]} | ({in2[21]} | ({in2[22]} | {in2[23]})));
 assign in1_31_0_ = ~(sub_407_2_n_34 & ~(sub_407_2_n_28 & {in1[38]}));
 assign sub_407_2_n_45 = ~({in2[12]} | ({in2[13]} | ({in2[14]} | {in2[15]})));
 assign sub_407_2_n_51 = ~(sub_407_2_n_41 | sub_407_2_n_1);
 assign sub_407_2_n_50 = ~(sub_407_2_n_4 | sub_407_2_n_35);
 assign sub_407_2_n_49 = ~(sub_407_2_n_9 | sub_407_2_n_35);
 assign sub_407_2_n_43 = ~sub_407_2_n_42;
 assign sub_407_2_n_44 = ~(in1_29_4_ & ~{in2[5]});
 assign sub_407_2_n_42 = ~(in1_29_3_ & ~{in2[4]});
 assign sub_407_2_n_41 = ~(sub_407_2_n_29 | ~sub_407_2_n_31);
 assign sub_407_2_n_40 = ~(sub_407_2_n_32 & {in2[3]});
 assign sub_407_2_n_39 = ~(in1_29_1_ & ~{in2[2]});
 assign sub_407_2_n_38 = ~(in1_29_1_ | ~{in2[2]});
 assign sub_407_2_n_25 = ~(in1_29_5_ & ~{in2[6]});
 assign sub_407_2_n_33 = ~(in1_29_0_ | sub_407_2_n_27);
 assign sub_407_2_n_37 = ~(in1_29_9_ & ~{in2[10]});
 assign sub_407_2_n_36 = ~(in1_29_7_ & ~{in2[8]});
 assign sub_407_2_n_35 = ~(in1_29_6_ | sub_407_2_n_30);
 assign sub_407_2_n_34 = ~({in2[0]} & ~{in1[38]});
 assign sub_407_2_n_32 = ~in1_29_2_;
 assign sub_407_2_n_31 = ~{in2[9]};
 assign sub_407_2_n_30 = ~{in2[7]};
 assign sub_407_2_n_29 = ~in1_29_8_;
 assign sub_407_2_n_28 = ~{in2[0]};
 assign sub_407_2_n_27 = ~{in2[1]};
 assign in1_31_2_ = ~(sub_407_2_n_14 ^ sub_407_2_n_74);
 assign in1_31_5_ = ~(sub_407_2_n_81 ^ sub_407_2_n_17);
 assign in1_31_3_ = (sub_407_2_n_80 ^ sub_407_2_n_15);
 assign in1_31_4_ = (sub_407_2_n_79 ^ sub_407_2_n_13);
 assign in1_31_6_ = ~(sub_407_2_n_82 ^ sub_407_2_n_12);
 assign sub_407_2_n_19 = ~(sub_407_2_n_78 | (sub_407_2_n_10 | ~sub_407_2_n_50));
 assign in1_31_7_ = (sub_407_2_n_84 ^ sub_407_2_n_49);
 assign sub_407_2_n_17 = ~(sub_407_2_n_3 | ~sub_407_2_n_44);
 assign sub_407_2_n_16 = (sub_407_2_n_37 & sub_407_2_n_8);
 assign sub_407_2_n_15 = (sub_407_2_n_40 & sub_407_2_n_7);
 assign sub_407_2_n_14 = ~(sub_407_2_n_38 | ~sub_407_2_n_39);
 assign sub_407_2_n_13 = ~(sub_407_2_n_43 | ~sub_407_2_n_2);
 assign sub_407_2_n_12 = ~(sub_407_2_n_4 | ~sub_407_2_n_25);
 assign sub_407_2_n_11 = ~(sub_407_2_n_6 | ~sub_407_2_n_36);
 assign sub_407_2_n_10 = ~(sub_407_2_n_2 & ~sub_407_2_n_3);
 assign sub_407_2_n_9 = (in1_29_6_ & sub_407_2_n_30);
 assign sub_407_2_n_8 = ~({in2[10]} & ~in1_29_9_);
 assign sub_407_2_n_7 = (sub_407_2_n_32 | {in2[3]});
 assign sub_407_2_n_6 = ~(in1_29_7_ | ~{in2[8]});
 assign sub_407_2_n_5 = ~(sub_407_2_n_8 & ~{in2[11]});
 assign sub_407_2_n_4 = ~(in1_29_5_ | ~{in2[6]});
 assign sub_407_2_n_3 = ~(in1_29_4_ | ~{in2[5]});
 assign sub_407_2_n_2 = ~({in2[4]} & ~in1_29_3_);
 assign sub_407_2_n_1 = ~(sub_407_2_n_31 | ~sub_407_2_n_29);
 assign sub_407_2_n_0 = (in1_29_0_ & sub_407_2_n_27);
 assign in1_34_11_ = ~((sub_426_2_n_68 & ~sub_426_2_n_120) | (sub_426_2_n_17 & sub_426_2_n_120));
 assign sub_426_2_n_120 = ~(sub_426_2_n_34 & (sub_426_2_n_22 | sub_426_2_n_30));
 assign in1_34_7_ = (sub_426_2_n_113 ^ sub_426_2_n_63);
 assign in1_34_9_ = ~(sub_426_2_n_116 & ~sub_426_2_n_117);
 assign sub_426_2_n_117 = ~(sub_426_2_n_112 | sub_426_2_n_62);
 assign sub_426_2_n_116 = ~(sub_426_2_n_112 & sub_426_2_n_62);
 assign in1_34_5_ = ~((sub_426_2_n_72 & ~sub_426_2_n_108) | (sub_426_2_n_12 & sub_426_2_n_108));
 assign in1_34_24_ = ~(sub_426_2_n_110 & sub_426_2_n_103);
 assign sub_426_2_n_113 = ~(sub_426_2_n_35 & (sub_426_2_n_105 | sub_426_2_n_4));
 assign sub_426_2_n_112 = ~(sub_426_2_n_51 | (sub_426_2_n_107 & sub_426_2_n_43));
 assign in1_34_8_ = ~((sub_426_2_n_54 & ~sub_426_2_n_107) | (sub_426_2_n_55 & sub_426_2_n_107));
 assign sub_426_2_n_110 = ~(sub_426_2_n_106 & sub_426_2_n_93);
 assign sub_426_2_n_109 = ~(sub_426_2_n_106 | sub_426_2_n_14);
 assign sub_426_2_n_108 = ~(sub_426_2_n_33 & (sub_426_2_n_101 | sub_426_2_n_5));
 assign sub_426_2_n_107 = ~sub_426_2_n_106;
 assign sub_426_2_n_106 = ~(sub_426_2_n_100 | sub_426_2_n_90);
 assign sub_426_2_n_105 = ~sub_426_2_n_104;
 assign sub_426_2_n_104 = ~(sub_426_2_n_80 & (sub_426_2_n_83 | sub_426_2_n_97));
 assign sub_426_2_n_103 = ~(sub_426_2_n_102 & sub_426_2_n_94);
 assign sub_426_2_n_102 = ~(sub_426_2_n_95 & (sub_426_2_n_75 | sub_426_2_n_1));
 assign sub_426_2_n_101 = ~(sub_426_2_n_96 | sub_426_2_n_76);
 assign sub_426_2_n_100 = (sub_426_2_n_98 & sub_426_2_n_85);
 assign sub_426_2_n_99 = ~(sub_426_2_n_91 & sub_426_2_n_50);
 assign sub_426_2_n_98 = ~(sub_426_2_n_91 & sub_426_2_n_67);
 assign sub_426_2_n_97 = (sub_426_2_n_11 & sub_426_2_n_67);
 assign sub_426_2_n_96 = ~(sub_426_2_n_11 | sub_426_2_n_66);
 assign sub_426_2_n_95 = (sub_426_2_n_23 & sub_426_2_n_42);
 assign sub_426_2_n_94 = ~(sub_426_2_n_77 & ~sub_426_2_n_89);
 assign sub_426_2_n_93 = ~(sub_426_2_n_84 | sub_426_2_n_77);
 assign in1_34_1_ = ~(in1_32_0_ ^ ({in2[1]} ^ sub_426_2_n_41));
 assign sub_426_2_n_91 = ~(sub_426_2_n_86 & sub_426_2_n_64);
 assign sub_426_2_n_90 = ~(sub_426_2_n_88 & sub_426_2_n_73);
 assign sub_426_2_n_89 = ~(sub_426_2_n_61 & (sub_426_2_n_58 & (sub_426_2_n_57 & sub_426_2_n_56)));
 assign sub_426_2_n_88 = ~(sub_426_2_n_79 & sub_426_2_n_71);
 assign sub_426_2_n_87 = ~(sub_426_2_n_2 | ~sub_426_2_n_41);
 assign sub_426_2_n_86 = ~(sub_426_2_n_46 & ~sub_426_2_n_41);
 assign sub_426_2_n_85 = ~(sub_426_2_n_82 | sub_426_2_n_10);
 assign sub_426_2_n_84 = ~(sub_426_2_n_74 | sub_426_2_n_9);
 assign sub_426_2_n_83 = ~(sub_426_2_n_78 & sub_426_2_n_81);
 assign sub_426_2_n_82 = ~(sub_426_2_n_70 & sub_426_2_n_49);
 assign sub_426_2_n_81 = ~(sub_426_2_n_67 & sub_426_2_n_7);
 assign sub_426_2_n_80 = ~sub_426_2_n_79;
 assign sub_426_2_n_79 = ~(sub_426_2_n_8 | (sub_426_2_n_33 & sub_426_2_n_47));
 assign sub_426_2_n_78 = (sub_426_2_n_65 & sub_426_2_n_70);
 assign sub_426_2_n_77 = ~(sub_426_2_n_53 & (sub_426_2_n_34 | sub_426_2_n_3));
 assign sub_426_2_n_76 = ~(sub_426_2_n_26 & (sub_426_2_n_50 | sub_426_2_n_29));
 assign sub_426_2_n_75 = ~(sub_426_2_n_31 | (sub_426_2_n_6 & sub_426_2_n_32));
 assign sub_426_2_n_74 = ~(sub_426_2_n_60 | sub_426_2_n_1);
 assign sub_426_2_n_73 = ~(sub_426_2_n_48 | ~(sub_426_2_n_35 | sub_426_2_n_45));
 assign sub_426_2_n_72 = ~sub_426_2_n_12;
 assign sub_426_2_n_71 = ~sub_426_2_n_10;
 assign sub_426_2_n_68 = ~sub_426_2_n_17;
 assign sub_426_2_n_66 = ~(sub_426_2_n_28 & ~sub_426_2_n_7);
 assign sub_426_2_n_65 = ~(sub_426_2_n_27 & sub_426_2_n_26);
 assign sub_426_2_n_64 = ~(sub_426_2_n_2 | sub_426_2_n_7);
 assign sub_426_2_n_63 = ~(sub_426_2_n_48 | sub_426_2_n_45);
 assign sub_426_2_n_70 = ~(sub_426_2_n_5 | sub_426_2_n_8);
 assign sub_426_2_n_69 = ~(sub_426_2_n_52 | sub_426_2_n_4);
 assign sub_426_2_n_67 = (sub_426_2_n_50 & sub_426_2_n_44);
 assign sub_426_2_n_61 = ~({in2[12]} | ({in2[13]} | {in2[14]}));
 assign sub_426_2_n_60 = ~(sub_426_2_n_32 | sub_426_2_n_31);
 assign in1_34_0_ = ~(sub_426_2_n_41 & ~(sub_426_2_n_38 & {in1[37]}));
 assign sub_426_2_n_58 = ~({in2[15]} | ({in2[16]} | {in2[17]}));
 assign sub_426_2_n_57 = ~({in2[18]} | ({in2[19]} | {in2[20]}));
 assign sub_426_2_n_56 = ~({in2[21]} | ({in2[22]} | {in2[23]}));
 assign sub_426_2_n_62 = ~(sub_426_2_n_1 | sub_426_2_n_31);
 assign sub_426_2_n_55 = ~(sub_426_2_n_51 | sub_426_2_n_6);
 assign sub_426_2_n_54 = ~(sub_426_2_n_32 & ~sub_426_2_n_6);
 assign sub_426_2_n_52 = ~sub_426_2_n_35;
 assign sub_426_2_n_51 = ~sub_426_2_n_32;
 assign sub_426_2_n_53 = ~(in1_32_10_ & ~{in2[11]});
 assign sub_426_2_n_35 = ~(sub_426_2_n_25 & ~{in2[6]});
 assign sub_426_2_n_34 = ~(in1_32_9_ & ~{in2[10]});
 assign sub_426_2_n_33 = ~(in1_32_3_ & ~{in2[4]});
 assign sub_426_2_n_32 = ~(in1_32_7_ & ~{in2[8]});
 assign sub_426_2_n_31 = ~(in1_32_8_ | sub_426_2_n_39);
 assign sub_426_2_n_50 = ~(in1_32_1_ & ~{in2[2]});
 assign sub_426_2_n_49 = (in1_32_2_ | sub_426_2_n_37);
 assign sub_426_2_n_43 = ~sub_426_2_n_6;
 assign sub_426_2_n_42 = ~sub_426_2_n_3;
 assign sub_426_2_n_48 = (sub_426_2_n_40 & in1_32_6_);
 assign sub_426_2_n_47 = ~(in1_32_4_ & ~{in2[5]});
 assign sub_426_2_n_46 = ~(in1_32_0_ & ~{in2[1]});
 assign sub_426_2_n_45 = ~(in1_32_6_ | sub_426_2_n_40);
 assign sub_426_2_n_30 = ~(in1_32_9_ | ~{in2[10]});
 assign sub_426_2_n_44 = ~(in1_32_2_ & ~{in2[3]});
 assign sub_426_2_n_41 = ~({in2[0]} & ~{in1[37]});
 assign sub_426_2_n_40 = ~{in2[7]};
 assign sub_426_2_n_39 = ~{in2[9]};
 assign sub_426_2_n_38 = ~{in2[0]};
 assign sub_426_2_n_37 = ~{in2[3]};
 assign sub_426_2_n_29 = ~sub_426_2_n_28;
 assign sub_426_2_n_28 = sub_426_2_n_49;
 assign sub_426_2_n_27 = ~sub_426_2_n_49;
 assign sub_426_2_n_26 = sub_426_2_n_44;
 assign sub_426_2_n_25 = in1_32_5_;
 assign in1_34_10_ = ~(sub_426_2_n_22 ^ sub_426_2_n_16);
 assign sub_426_2_n_23 = ~(sub_426_2_n_30 | sub_426_2_n_89);
 assign sub_426_2_n_22 = ~(sub_426_2_n_109 | ~sub_426_2_n_74);
 assign in1_34_6_ = (sub_426_2_n_104 ^ sub_426_2_n_69);
 assign in1_34_3_ = (sub_426_2_n_99 ^ sub_426_2_n_0);
 assign in1_34_2_ = ~(sub_426_2_n_11 ^ sub_426_2_n_13);
 assign in1_34_4_ = ~(sub_426_2_n_101 ^ sub_426_2_n_15);
 assign sub_426_2_n_17 = ~(sub_426_2_n_3 | ~sub_426_2_n_53);
 assign sub_426_2_n_16 = ~(sub_426_2_n_30 | ~sub_426_2_n_34);
 assign sub_426_2_n_15 = ~(sub_426_2_n_5 | ~sub_426_2_n_33);
 assign sub_426_2_n_14 = ~(sub_426_2_n_43 & ~sub_426_2_n_31);
 assign sub_426_2_n_13 = ~(sub_426_2_n_7 | ~sub_426_2_n_50);
 assign sub_426_2_n_12 = ~(sub_426_2_n_8 | ~sub_426_2_n_47);
 assign sub_426_2_n_11 = ~(sub_426_2_n_87 | ~sub_426_2_n_46);
 assign sub_426_2_n_10 = (sub_426_2_n_45 | sub_426_2_n_4);
 assign sub_426_2_n_9 = ~(sub_426_2_n_42 & ~sub_426_2_n_30);
 assign sub_426_2_n_8 = ~(in1_32_4_ | ~{in2[5]});
 assign sub_426_2_n_7 = ~(in1_32_1_ | ~{in2[2]});
 assign sub_426_2_n_6 = ~(in1_32_7_ | ~{in2[8]});
 assign sub_426_2_n_5 = ~(in1_32_3_ | ~{in2[4]});
 assign sub_426_2_n_4 = ~(in1_32_5_ | ~{in2[6]});
 assign sub_426_2_n_3 = ~(in1_32_10_ | ~{in2[11]});
 assign sub_426_2_n_2 = ~(in1_32_0_ | ~{in2[1]});
 assign sub_426_2_n_1 = (in1_32_8_ & sub_426_2_n_39);
 assign sub_426_2_n_0 = ~(sub_426_2_n_29 | ~sub_426_2_n_26);
 assign in1_37_11_ = (sub_445_2_n_143 ^ sub_445_2_n_69);
 assign in1_37_9_ = ~((sub_445_2_n_77 & ~sub_445_2_n_138) | (sub_445_2_n_76 & sub_445_2_n_138));
 assign in1_37_12_ = (sub_445_2_n_136 ^ sub_445_2_n_59);
 assign sub_445_2_n_143 = ~(sub_445_2_n_55 & (sub_445_2_n_133 | sub_445_2_n_56));
 assign in1_37_10_ = ~(sub_445_2_n_141 & ~sub_445_2_n_140);
 assign sub_445_2_n_141 = ~(sub_445_2_n_134 & sub_445_2_n_78);
 assign sub_445_2_n_140 = ~(sub_445_2_n_134 | sub_445_2_n_78);
 assign in1_37_24_ = ~(sub_445_2_n_128 & sub_445_2_n_131);
 assign sub_445_2_n_138 = ~(sub_445_2_n_42 & (sub_445_2_n_126 | sub_445_2_n_2));
 assign sub_445_2_n_137 = ~(sub_445_2_n_45 & (sub_445_2_n_129 | sub_445_2_n_43));
 assign sub_445_2_n_136 = ~(sub_445_2_n_25 & (sub_445_2_n_126 | sub_445_2_n_17));
 assign in1_37_8_ = ~(sub_445_2_n_126 ^ sub_445_2_n_12);
 assign sub_445_2_n_134 = ~sub_445_2_n_133;
 assign sub_445_2_n_133 = ~(sub_445_2_n_109 | sub_445_2_n_130);
 assign sub_445_2_n_132 = ~(sub_445_2_n_57 & (sub_445_2_n_120 | sub_445_2_n_28));
 assign sub_445_2_n_131 = ~(sub_445_2_n_127 & sub_445_2_n_25);
 assign sub_445_2_n_130 = ~(sub_445_2_n_118 | sub_445_2_n_29);
 assign sub_445_2_n_129 = ~(sub_445_2_n_87 | (sub_445_2_n_95 & sub_445_2_n_112));
 assign sub_445_2_n_128 = ~(sub_445_2_n_121 & sub_445_2_n_117);
 assign sub_445_2_n_127 = ~(sub_445_2_n_122 | sub_445_2_n_101);
 assign sub_445_2_n_126 = ~(sub_445_2_n_119 | sub_445_2_n_24);
 assign in1_37_3_ = ~(sub_445_2_n_124 & ~sub_445_2_n_123);
 assign sub_445_2_n_124 = ~(sub_445_2_n_116 & sub_445_2_n_79);
 assign sub_445_2_n_123 = ~(sub_445_2_n_116 | sub_445_2_n_79);
 assign sub_445_2_n_122 = ~(sub_445_2_n_107 | sub_445_2_n_111);
 assign sub_445_2_n_121 = ~(sub_445_2_n_114 | sub_445_2_n_26);
 assign sub_445_2_n_120 = ~(sub_445_2_n_110 | sub_445_2_n_83);
 assign sub_445_2_n_119 = ~sub_445_2_n_118;
 assign sub_445_2_n_118 = ~(sub_445_2_n_113 & sub_445_2_n_94);
 assign sub_445_2_n_117 = ~(sub_445_2_n_115 & sub_445_2_n_98);
 assign sub_445_2_n_116 = ~(sub_445_2_n_103 & sub_445_2_n_53);
 assign sub_445_2_n_115 = ~(sub_445_2_n_105 | sub_445_2_n_14);
 assign sub_445_2_n_114 = ~(sub_445_2_n_105 | sub_445_2_n_86);
 assign sub_445_2_n_113 = ~(sub_445_2_n_103 & sub_445_2_n_32);
 assign sub_445_2_n_112 = ~(sub_445_2_n_11 & sub_445_2_n_32);
 assign sub_445_2_n_111 = ~(sub_445_2_n_89 | ~sub_445_2_n_103);
 assign sub_445_2_n_110 = ~(sub_445_2_n_11 | sub_445_2_n_71);
 assign sub_445_2_n_109 = ~(sub_445_2_n_106 & sub_445_2_n_108);
 assign sub_445_2_n_108 = ~(sub_445_2_n_92 & sub_445_2_n_30);
 assign sub_445_2_n_107 = ~(sub_445_2_n_93 & sub_445_2_n_88);
 assign sub_445_2_n_106 = (sub_445_2_n_100 & sub_445_2_n_84);
 assign sub_445_2_n_105 = ~(sub_445_2_n_102 & (in1_35_11_ | sub_445_2_n_36));
 assign in1_37_1_ = ~(in1_35_0_ ^ ({in2[1]} ^ sub_445_2_n_51));
 assign sub_445_2_n_103 = ~(sub_445_2_n_96 & sub_445_2_n_65);
 assign sub_445_2_n_102 = ~(sub_445_2_n_90 | ~sub_445_2_n_68);
 assign sub_445_2_n_101 = ~(sub_445_2_n_19 & ~sub_445_2_n_85);
 assign sub_445_2_n_100 = ~(sub_445_2_n_85 & sub_445_2_n_30);
 assign sub_445_2_n_99 = ~(sub_445_2_n_44 | ~sub_445_2_n_51);
 assign sub_445_2_n_98 = ~(sub_445_2_n_84 & sub_445_2_n_29);
 assign sub_445_2_n_97 = ~(sub_445_2_n_84 | sub_445_2_n_14);
 assign sub_445_2_n_96 = ~(sub_445_2_n_41 & ~sub_445_2_n_51);
 assign sub_445_2_n_95 = ~(sub_445_2_n_81 | sub_445_2_n_20);
 assign sub_445_2_n_94 = (sub_445_2_n_82 & sub_445_2_n_73);
 assign sub_445_2_n_93 = ~(sub_445_2_n_80 | sub_445_2_n_74);
 assign sub_445_2_n_92 = ~(sub_445_2_n_31 | (sub_445_2_n_74 | ~sub_445_2_n_7));
 assign sub_445_2_n_91 = ~(sub_445_2_n_67 & (sub_445_2_n_73 & ~sub_445_2_n_40));
 assign sub_445_2_n_89 = ~(sub_445_2_n_32 & sub_445_2_n_31);
 assign sub_445_2_n_88 = ~(sub_445_2_n_31 & ~sub_445_2_n_39);
 assign sub_445_2_n_87 = ~(sub_445_2_n_31 | sub_445_2_n_40);
 assign sub_445_2_n_90 = ~(sub_445_2_n_64 & sub_445_2_n_63);
 assign sub_445_2_n_83 = ~(sub_445_2_n_52 & (sub_445_2_n_53 | sub_445_2_n_4));
 assign sub_445_2_n_82 = ~(sub_445_2_n_28 | (sub_445_2_n_40 | sub_445_2_n_4));
 assign sub_445_2_n_81 = ~(sub_445_2_n_70 & sub_445_2_n_60);
 assign sub_445_2_n_80 = ~(sub_445_2_n_7 & ~(sub_445_2_n_28 & sub_445_2_n_48));
 assign sub_445_2_n_86 = ~(sub_445_2_n_72 | sub_445_2_n_9);
 assign sub_445_2_n_85 = ~(sub_445_2_n_58 & (sub_445_2_n_45 | sub_445_2_n_0));
 assign sub_445_2_n_84 = ~(sub_445_2_n_66 | sub_445_2_n_10);
 assign sub_445_2_n_77 = ~sub_445_2_n_76;
 assign sub_445_2_n_73 = ~sub_445_2_n_74;
 assign sub_445_2_n_72 = ~(sub_445_2_n_55 | sub_445_2_n_46);
 assign sub_445_2_n_71 = ~(sub_445_2_n_39 & ~sub_445_2_n_3);
 assign sub_445_2_n_70 = ~(sub_445_2_n_4 & sub_445_2_n_52);
 assign sub_445_2_n_79 = ~(sub_445_2_n_52 & sub_445_2_n_39);
 assign sub_445_2_n_78 = ~(sub_445_2_n_55 & sub_445_2_n_6);
 assign sub_445_2_n_76 = ~(sub_445_2_n_10 | sub_445_2_n_47);
 assign sub_445_2_n_69 = ~(sub_445_2_n_9 | sub_445_2_n_46);
 assign sub_445_2_n_75 = ~(sub_445_2_n_49 | sub_445_2_n_40);
 assign sub_445_2_n_74 = ~(sub_445_2_n_8 & sub_445_2_n_54);
 assign sub_445_2_n_32 = (sub_445_2_n_53 & sub_445_2_n_52);
 assign sub_445_2_n_67 = ~sub_445_2_n_31;
 assign sub_445_2_n_29 = ~sub_445_2_n_30;
 assign sub_445_2_n_66 = ~(sub_445_2_n_42 | sub_445_2_n_47);
 assign sub_445_2_n_65 = ~(sub_445_2_n_44 | sub_445_2_n_3);
 assign sub_445_2_n_64 = ~({in2[16]} | ({in2[17]} | ({in2[18]} | {in2[19]})));
 assign sub_445_2_n_63 = ~({in2[20]} | ({in2[21]} | ({in2[22]} | {in2[23]})));
 assign in1_37_0_ = ~(sub_445_2_n_51 & ~(sub_445_2_n_37 & {in1[36]}));
 assign sub_445_2_n_61 = ~(sub_445_2_n_1 | sub_445_2_n_28);
 assign sub_445_2_n_60 = ~(sub_445_2_n_28 | sub_445_2_n_40);
 assign sub_445_2_n_68 = ~({in2[14]} | ({in2[15]} | {in2[13]}));
 assign sub_445_2_n_59 = ~(sub_445_2_n_5 | sub_445_2_n_50);
 assign sub_445_2_n_31 = ~(sub_445_2_n_1 | sub_445_2_n_49);
 assign sub_445_2_n_30 = ~(sub_445_2_n_2 | sub_445_2_n_47);
 assign sub_445_2_n_57 = ~sub_445_2_n_1;
 assign sub_445_2_n_56 = ~sub_445_2_n_6;
 assign sub_445_2_n_54 = ~sub_445_2_n_0;
 assign sub_445_2_n_58 = ~(in1_35_6_ & ~{in2[7]});
 assign sub_445_2_n_50 = ~(in1_35_11_ | sub_445_2_n_36);
 assign sub_445_2_n_55 = ~(in1_35_9_ & ~{in2[10]});
 assign sub_445_2_n_53 = ~(in1_35_1_ & ~{in2[2]});
 assign sub_445_2_n_52 = ~(in1_35_2_ & ~{in2[3]});
 assign sub_445_2_n_51 = ~({in2[0]} & ~{in1[36]});
 assign sub_445_2_n_49 = ~sub_445_2_n_48;
 assign sub_445_2_n_43 = ~sub_445_2_n_8;
 assign sub_445_2_n_40 = ~sub_445_2_n_7;
 assign sub_445_2_n_39 = ~sub_445_2_n_4;
 assign sub_445_2_n_48 = ~(in1_35_4_ & ~{in2[5]});
 assign sub_445_2_n_47 = ~(in1_35_8_ | sub_445_2_n_35);
 assign sub_445_2_n_46 = ~(in1_35_10_ | sub_445_2_n_34);
 assign sub_445_2_n_45 = ~(in1_35_5_ & ~{in2[6]});
 assign sub_445_2_n_44 = ~(in1_35_0_ | ~{in2[1]});
 assign sub_445_2_n_42 = ~(in1_35_7_ & ~{in2[8]});
 assign sub_445_2_n_41 = ~(in1_35_0_ & ~{in2[1]});
 assign sub_445_2_n_38 = ~{in2[4]};
 assign sub_445_2_n_37 = ~{in2[0]};
 assign sub_445_2_n_36 = ~{in2[12]};
 assign sub_445_2_n_35 = ~{in2[9]};
 assign sub_445_2_n_34 = ~{in2[11]};
 assign sub_445_2_n_28 = ~(in1_35_3_ | sub_445_2_n_38);
 assign in1_37_4_ = ~(sub_445_2_n_120 ^ sub_445_2_n_61);
 assign sub_445_2_n_26 = ~(sub_445_2_n_19 | sub_445_2_n_90);
 assign sub_445_2_n_25 = ~(sub_445_2_n_97 | ~sub_445_2_n_86);
 assign sub_445_2_n_24 = ~(sub_445_2_n_91 & ~sub_445_2_n_85);
 assign in1_37_6_ = ~(sub_445_2_n_129 ^ sub_445_2_n_13);
 assign in1_37_7_ = (sub_445_2_n_137 ^ sub_445_2_n_16);
 assign in1_37_5_ = (sub_445_2_n_132 ^ sub_445_2_n_75);
 assign sub_445_2_n_20 = (sub_445_2_n_32 & sub_445_2_n_3);
 assign sub_445_2_n_19 = ~(sub_445_2_n_5 & sub_445_2_n_68);
 assign in1_37_2_ = ~(sub_445_2_n_11 ^ sub_445_2_n_15);
 assign sub_445_2_n_17 = ~(sub_445_2_n_30 & ~sub_445_2_n_14);
 assign sub_445_2_n_16 = ~(sub_445_2_n_0 | ~sub_445_2_n_58);
 assign sub_445_2_n_15 = ~(sub_445_2_n_3 | ~sub_445_2_n_53);
 assign sub_445_2_n_14 = ~(sub_445_2_n_6 & ~sub_445_2_n_46);
 assign sub_445_2_n_13 = ~(sub_445_2_n_43 | ~sub_445_2_n_45);
 assign sub_445_2_n_12 = ~(sub_445_2_n_2 | ~sub_445_2_n_42);
 assign sub_445_2_n_11 = ~(sub_445_2_n_99 | ~sub_445_2_n_41);
 assign sub_445_2_n_10 = (in1_35_8_ & sub_445_2_n_35);
 assign sub_445_2_n_9 = (in1_35_10_ & sub_445_2_n_34);
 assign sub_445_2_n_8 = ~({in2[6]} & ~in1_35_5_);
 assign sub_445_2_n_7 = ~({in2[5]} & ~in1_35_4_);
 assign sub_445_2_n_6 = ~({in2[10]} & ~in1_35_9_);
 assign sub_445_2_n_5 = (in1_35_11_ & sub_445_2_n_36);
 assign sub_445_2_n_4 = ~(in1_35_2_ | ~{in2[3]});
 assign sub_445_2_n_3 = ~(in1_35_1_ | ~{in2[2]});
 assign sub_445_2_n_2 = ~(in1_35_7_ | ~{in2[8]});
 assign sub_445_2_n_1 = (in1_35_3_ & sub_445_2_n_38);
 assign sub_445_2_n_0 = ~(in1_35_6_ | ~{in2[7]});
 assign in1_40_13_ = (sub_466_2_n_147 ^ sub_466_2_n_68);
 assign sub_466_2_n_147 = ~(sub_466_2_n_50 & (sub_466_2_n_137 | sub_466_2_n_35));
 assign sub_466_2_n_146 = ~(sub_466_2_n_62 & (sub_466_2_n_139 | sub_466_2_n_1));
 assign in1_40_10_ = ~(sub_466_2_n_139 ^ sub_466_2_n_17);
 assign sub_466_2_n_144 = ~(sub_466_2_n_65 & (sub_466_2_n_135 | sub_466_2_n_53));
 assign in1_40_6_ = ~(sub_466_2_n_140 & ~sub_466_2_n_141);
 assign in1_40_24_ = ~(sub_466_2_n_95 & (sub_466_2_n_134 | sub_466_2_n_125));
 assign sub_466_2_n_141 = ~(sub_466_2_n_135 | sub_466_2_n_18);
 assign sub_466_2_n_140 = ~(sub_466_2_n_135 & sub_466_2_n_18);
 assign sub_466_2_n_139 = ~(sub_466_2_n_116 | sub_466_2_n_26);
 assign sub_466_2_n_138 = ~(sub_466_2_n_67 & (sub_466_2_n_130 | sub_466_2_n_54));
 assign sub_466_2_n_137 = ~(sub_466_2_n_136 | sub_466_2_n_114);
 assign sub_466_2_n_136 = ~(sub_466_2_n_130 | sub_466_2_n_97);
 assign sub_466_2_n_135 = ~(sub_466_2_n_92 | (sub_466_2_n_39 & sub_466_2_n_33));
 assign sub_466_2_n_134 = ~(sub_466_2_n_131 | sub_466_2_n_119);
 assign sub_466_2_n_133 = ~(sub_466_2_n_55 & (sub_466_2_n_123 | sub_466_2_n_34));
 assign in1_40_3_ = ~(sub_466_2_n_129 & ~sub_466_2_n_128);
 assign sub_466_2_n_131 = ~(sub_466_2_n_127 & sub_466_2_n_111);
 assign sub_466_2_n_130 = ~(sub_466_2_n_126 | sub_466_2_n_110);
 assign sub_466_2_n_129 = ~(sub_466_2_n_120 & sub_466_2_n_86);
 assign sub_466_2_n_128 = ~(sub_466_2_n_120 | sub_466_2_n_86);
 assign sub_466_2_n_127 = ~(sub_466_2_n_117 & sub_466_2_n_99);
 assign sub_466_2_n_126 = ~(sub_466_2_n_117 | sub_466_2_n_108);
 assign sub_466_2_n_125 = ~(sub_466_2_n_118 | sub_466_2_n_21);
 assign in1_40_2_ = ~(sub_466_2_n_121 & ~sub_466_2_n_122);
 assign sub_466_2_n_123 = ~sub_466_2_n_39;
 assign sub_466_2_n_39 = ~(sub_466_2_n_15 & (sub_466_2_n_113 | sub_466_2_n_73));
 assign sub_466_2_n_122 = ~(sub_466_2_n_113 | sub_466_2_n_14);
 assign sub_466_2_n_121 = ~(sub_466_2_n_113 & sub_466_2_n_14);
 assign sub_466_2_n_120 = ~(sub_466_2_n_31 & sub_466_2_n_59);
 assign sub_466_2_n_119 = ~(sub_466_2_n_89 & (sub_466_2_n_106 | sub_466_2_n_38));
 assign sub_466_2_n_118 = ~(sub_466_2_n_115 & sub_466_2_n_107);
 assign sub_466_2_n_117 = ~(sub_466_2_n_23 & sub_466_2_n_94);
 assign sub_466_2_n_116 = ~(sub_466_2_n_112 & sub_466_2_n_104);
 assign sub_466_2_n_115 = ~(sub_466_2_n_102 & sub_466_2_n_74);
 assign sub_466_2_n_114 = ~(sub_466_2_n_102 | sub_466_2_n_98);
 assign sub_466_2_n_113 = ~(sub_466_2_n_105 | sub_466_2_n_8);
 assign sub_466_2_n_112 = ~(sub_466_2_n_93 | (sub_466_2_n_38 & sub_466_2_n_82));
 assign sub_466_2_n_111 = ~(sub_466_2_n_103 | sub_466_2_n_97);
 assign sub_466_2_n_110 = ~(sub_466_2_n_37 & (sub_466_2_n_91 | sub_466_2_n_16));
 assign in1_40_1_ = ~(sub_466_2_n_101 & ~sub_466_2_n_100);
 assign sub_466_2_n_108 = (sub_466_2_n_96 | sub_466_2_n_16);
 assign sub_466_2_n_107 = ~(sub_466_2_n_98 & sub_466_2_n_74);
 assign sub_466_2_n_106 = ~(sub_466_2_n_96 & sub_466_2_n_91);
 assign sub_466_2_n_105 = ~(sub_466_2_n_61 | ~sub_466_2_n_49);
 assign sub_466_2_n_104 = ~(sub_466_2_n_92 & ~sub_466_2_n_20);
 assign sub_466_2_n_103 = ~(sub_466_2_n_38 | ~sub_466_2_n_16);
 assign sub_466_2_n_101 = ~(sub_466_2_n_88 & sub_466_2_n_49);
 assign sub_466_2_n_100 = ~(sub_466_2_n_88 | sub_466_2_n_49);
 assign sub_466_2_n_99 = (sub_466_2_n_91 & sub_466_2_n_37);
 assign sub_466_2_n_102 = ~(sub_466_2_n_93 | sub_466_2_n_70);
 assign sub_466_2_n_95 = (sub_466_2_n_71 & sub_466_2_n_72);
 assign sub_466_2_n_94 = (sub_466_2_n_33 & sub_466_2_n_4);
 assign sub_466_2_n_98 = ~(sub_466_2_n_84 | sub_466_2_n_64);
 assign sub_466_2_n_97 = ~(sub_466_2_n_82 & sub_466_2_n_84);
 assign sub_466_2_n_96 = ~(sub_466_2_n_76 | sub_466_2_n_83);
 assign sub_466_2_n_38 = ~sub_466_2_n_37;
 assign sub_466_2_n_92 = ~sub_466_2_n_91;
 assign sub_466_2_n_90 = ~(sub_466_2_n_58 | (sub_466_2_n_57 & sub_466_2_n_51));
 assign sub_466_2_n_89 = ~(sub_466_2_n_81 | sub_466_2_n_35);
 assign sub_466_2_n_93 = ~(sub_466_2_n_66 & (sub_466_2_n_48 | sub_466_2_n_5));
 assign sub_466_2_n_37 = ~(sub_466_2_n_80 | sub_466_2_n_11);
 assign sub_466_2_n_91 = ~(sub_466_2_n_79 | sub_466_2_n_2);
 assign sub_466_2_n_81 = ~(sub_466_2_n_9 & ~sub_466_2_n_58);
 assign sub_466_2_n_80 = ~(sub_466_2_n_65 | sub_466_2_n_36);
 assign sub_466_2_n_79 = ~(sub_466_2_n_55 | sub_466_2_n_56);
 assign sub_466_2_n_88 = (sub_466_2_n_8 | sub_466_2_n_61);
 assign sub_466_2_n_87 = ~(sub_466_2_n_64 | sub_466_2_n_10);
 assign sub_466_2_n_86 = ~(sub_466_2_n_60 & sub_466_2_n_4);
 assign sub_466_2_n_78 = ~(sub_466_2_n_6 | sub_466_2_n_35);
 assign sub_466_2_n_85 = ~(sub_466_2_n_7 | sub_466_2_n_54);
 assign sub_466_2_n_84 = ~(sub_466_2_n_1 | sub_466_2_n_10);
 assign sub_466_2_n_83 = ~(sub_466_2_n_61 | sub_466_2_n_0);
 assign sub_466_2_n_82 = ~(sub_466_2_n_54 | sub_466_2_n_5);
 assign sub_466_2_n_73 = ~(sub_466_2_n_4 & ~sub_466_2_n_0);
 assign sub_466_2_n_72 = ~({in2[20]} | ({in2[21]} | ({in2[22]} | {in2[23]})));
 assign sub_466_2_n_71 = ~({in2[16]} | ({in2[17]} | ({in2[18]} | {in2[19]})));
 assign sub_466_2_n_70 = ~(sub_466_2_n_62 & sub_466_2_n_63);
 assign in1_40_0_ = ~(sub_466_2_n_49 & ~(sub_466_2_n_46 & {in1[35]}));
 assign sub_466_2_n_77 = ~(sub_466_2_n_11 | sub_466_2_n_36);
 assign sub_466_2_n_76 = ~(sub_466_2_n_59 & sub_466_2_n_60);
 assign sub_466_2_n_68 = ~(sub_466_2_n_52 | sub_466_2_n_57);
 assign sub_466_2_n_75 = ~(sub_466_2_n_2 | sub_466_2_n_56);
 assign sub_466_2_n_74 = ~(sub_466_2_n_6 | sub_466_2_n_52);
 assign sub_466_2_n_67 = ~sub_466_2_n_7;
 assign sub_466_2_n_64 = ~sub_466_2_n_63;
 assign sub_466_2_n_66 = ~(in1_38_8_ & ~{in2[9]});
 assign sub_466_2_n_65 = ~(in1_38_5_ & ~{in2[6]});
 assign sub_466_2_n_63 = ~(in1_38_10_ & ~{in2[11]});
 assign sub_466_2_n_62 = ~(in1_38_9_ & ~{in2[10]});
 assign sub_466_2_n_61 = ~(in1_38_0_ | sub_466_2_n_42);
 assign sub_466_2_n_36 = ~(in1_38_6_ | sub_466_2_n_44);
 assign sub_466_2_n_60 = ~(in1_38_2_ & ~{in2[3]});
 assign sub_466_2_n_59 = ~(in1_38_1_ & ~{in2[2]});
 assign sub_466_2_n_57 = ~sub_466_2_n_9;
 assign sub_466_2_n_53 = ~sub_466_2_n_3;
 assign sub_466_2_n_52 = ~sub_466_2_n_51;
 assign sub_466_2_n_50 = ~sub_466_2_n_6;
 assign sub_466_2_n_48 = ~(in1_38_7_ & ~{in2[8]});
 assign sub_466_2_n_58 = ({in2[14]} | {in2[15]});
 assign sub_466_2_n_56 = ~(in1_38_4_ | sub_466_2_n_43);
 assign sub_466_2_n_55 = ~(in1_38_3_ & ~{in2[4]});
 assign sub_466_2_n_54 = ~(in1_38_7_ | sub_466_2_n_41);
 assign sub_466_2_n_51 = ~(in1_38_12_ & ~{in2[13]});
 assign sub_466_2_n_35 = ~(in1_38_11_ | sub_466_2_n_45);
 assign sub_466_2_n_49 = ~({in2[0]} & ~{in1[35]});
 assign sub_466_2_n_47 = ~{in2[4]};
 assign sub_466_2_n_46 = ~{in2[0]};
 assign sub_466_2_n_45 = ~{in2[12]};
 assign sub_466_2_n_44 = ~{in2[7]};
 assign sub_466_2_n_43 = ~{in2[5]};
 assign sub_466_2_n_42 = ~{in2[1]};
 assign sub_466_2_n_41 = ~{in2[8]};
 assign sub_466_2_n_34 = ~(in1_38_3_ | sub_466_2_n_47);
 assign sub_466_2_n_33 = ~(sub_466_2_n_34 | sub_466_2_n_56);
 assign in1_40_12_ = ~(sub_466_2_n_137 ^ sub_466_2_n_78);
 assign sub_466_2_n_31 = ~(sub_466_2_n_83 & ~sub_466_2_n_30);
 assign sub_466_2_n_30 = ~(sub_466_2_n_8 | sub_466_2_n_49);
 assign in1_40_11_ = (sub_466_2_n_146 ^ sub_466_2_n_87);
 assign in1_40_8_ = ~(sub_466_2_n_130 ^ sub_466_2_n_85);
 assign in1_40_9_ = (sub_466_2_n_138 ^ sub_466_2_n_19);
 assign sub_466_2_n_26 = ~(sub_466_2_n_123 | (sub_466_2_n_20 | ~sub_466_2_n_33));
 assign in1_40_4_ = (sub_466_2_n_39 ^ sub_466_2_n_13);
 assign in1_40_7_ = (sub_466_2_n_144 ^ sub_466_2_n_77);
 assign sub_466_2_n_23 = ~(sub_466_2_n_30 & ~sub_466_2_n_76);
 assign in1_40_5_ = (sub_466_2_n_133 ^ sub_466_2_n_75);
 assign sub_466_2_n_21 = ~(sub_466_2_n_90 & ~(sub_466_2_n_74 & sub_466_2_n_35));
 assign sub_466_2_n_20 = ~(sub_466_2_n_82 & ~sub_466_2_n_16);
 assign sub_466_2_n_19 = ~(sub_466_2_n_5 | ~sub_466_2_n_66);
 assign sub_466_2_n_18 = ~(sub_466_2_n_53 | ~sub_466_2_n_65);
 assign sub_466_2_n_17 = ~(sub_466_2_n_1 | ~sub_466_2_n_62);
 assign sub_466_2_n_16 = ~(sub_466_2_n_3 & ~sub_466_2_n_36);
 assign sub_466_2_n_15 = ~(sub_466_2_n_12 | ~sub_466_2_n_60);
 assign sub_466_2_n_14 = ~(sub_466_2_n_0 | ~sub_466_2_n_59);
 assign sub_466_2_n_13 = ~(sub_466_2_n_34 | ~sub_466_2_n_55);
 assign sub_466_2_n_12 = ~(sub_466_2_n_59 | ~sub_466_2_n_4);
 assign sub_466_2_n_11 = (in1_38_6_ & sub_466_2_n_44);
 assign sub_466_2_n_10 = ~(in1_38_10_ | ~{in2[11]});
 assign sub_466_2_n_9 = ~({in2[13]} & ~in1_38_12_);
 assign sub_466_2_n_8 = (in1_38_0_ & sub_466_2_n_42);
 assign sub_466_2_n_7 = (in1_38_7_ & sub_466_2_n_41);
 assign sub_466_2_n_6 = (in1_38_11_ & sub_466_2_n_45);
 assign sub_466_2_n_5 = ~(in1_38_8_ | ~{in2[9]});
 assign sub_466_2_n_4 = ~({in2[3]} & ~in1_38_2_);
 assign sub_466_2_n_3 = ~({in2[6]} & ~in1_38_5_);
 assign sub_466_2_n_2 = (in1_38_4_ & sub_466_2_n_43);
 assign sub_466_2_n_1 = ~(in1_38_9_ | ~{in2[10]});
 assign sub_466_2_n_0 = ~(in1_38_1_ | ~{in2[2]});
 assign in1_43_14_ = (sub_487_2_n_127 ^ sub_487_2_n_20);
 assign in1_43_13_ = (sub_487_2_n_126 ^ sub_487_2_n_24);
 assign in1_43_11_ = (sub_487_2_n_125 ^ sub_487_2_n_71);
 assign in1_43_24_ = ~(sub_487_2_n_124 & sub_487_2_n_91);
 assign sub_487_2_n_127 = ~(sub_487_2_n_87 & (sub_487_2_n_34 | sub_487_2_n_80));
 assign sub_487_2_n_126 = ~(sub_487_2_n_38 & (sub_487_2_n_34 | sub_487_2_n_1));
 assign sub_487_2_n_125 = ~(sub_487_2_n_44 & (sub_487_2_n_118 | sub_487_2_n_6));
 assign sub_487_2_n_124 = ~(sub_487_2_n_123 & sub_487_2_n_110);
 assign sub_487_2_n_123 = ~(sub_487_2_n_119 & sub_487_2_n_94);
 assign sub_487_2_n_122 = ~(sub_487_2_n_43 & (sub_487_2_n_117 | sub_487_2_n_5));
 assign sub_487_2_n_121 = ~(sub_487_2_n_49 & (sub_487_2_n_116 | sub_487_2_n_8));
 assign in1_43_6_ = ~(sub_487_2_n_115 ^ sub_487_2_n_70);
 assign sub_487_2_n_119 = ~(sub_487_2_n_117 | sub_487_2_n_92);
 assign sub_487_2_n_118 = ~(sub_487_2_n_113 | (sub_487_2_n_35 | ~sub_487_2_n_88));
 assign sub_487_2_n_117 = ~(sub_487_2_n_112 | sub_487_2_n_102);
 assign sub_487_2_n_116 = ~sub_487_2_n_115;
 assign sub_487_2_n_115 = ~(sub_487_2_n_22 & (sub_487_2_n_109 | sub_487_2_n_65));
 assign sub_487_2_n_114 = ~(sub_487_2_n_37 & (sub_487_2_n_109 | sub_487_2_n_11));
 assign sub_487_2_n_113 = ~(sub_487_2_n_95 | sub_487_2_n_111);
 assign sub_487_2_n_112 = ~(sub_487_2_n_111 | sub_487_2_n_96);
 assign sub_487_2_n_111 = ~(sub_487_2_n_107 | sub_487_2_n_14);
 assign sub_487_2_n_110 = ~(sub_487_2_n_108 | sub_487_2_n_105);
 assign sub_487_2_n_109 = ~(sub_487_2_n_106 | sub_487_2_n_83);
 assign sub_487_2_n_108 = ~(sub_487_2_n_101 | ~sub_487_2_n_94);
 assign sub_487_2_n_107 = ~(sub_487_2_n_103 & sub_487_2_n_47);
 assign sub_487_2_n_106 = ~(sub_487_2_n_17 | sub_487_2_n_63);
 assign sub_487_2_n_105 = ~(sub_487_2_n_72 & ~(sub_487_2_n_86 & sub_487_2_n_82));
 assign in1_43_1_ = ~(sub_487_2_n_99 & ~sub_487_2_n_98);
 assign sub_487_2_n_103 = ~(sub_487_2_n_97 & sub_487_2_n_62);
 assign sub_487_2_n_102 = ~(sub_487_2_n_89 & (sub_487_2_n_22 | sub_487_2_n_78));
 assign sub_487_2_n_101 = ~(sub_487_2_n_29 | sub_487_2_n_84);
 assign sub_487_2_n_100 = ~(sub_487_2_n_7 | ~sub_487_2_n_53);
 assign sub_487_2_n_99 = ~(sub_487_2_n_66 & sub_487_2_n_53);
 assign sub_487_2_n_98 = ~(sub_487_2_n_66 | sub_487_2_n_53);
 assign sub_487_2_n_97 = ~(sub_487_2_n_45 & ~sub_487_2_n_53);
 assign sub_487_2_n_96 = ~(sub_487_2_n_90 & sub_487_2_n_64);
 assign sub_487_2_n_95 = ~(sub_487_2_n_85 & sub_487_2_n_93);
 assign sub_487_2_n_93 = ~(sub_487_2_n_65 | sub_487_2_n_78);
 assign sub_487_2_n_92 = ~(sub_487_2_n_75 & sub_487_2_n_69);
 assign sub_487_2_n_91 = (sub_487_2_n_58 & sub_487_2_n_61);
 assign sub_487_2_n_90 = (sub_487_2_n_77 & sub_487_2_n_9);
 assign sub_487_2_n_89 = ~(sub_487_2_n_73 | sub_487_2_n_12);
 assign sub_487_2_n_94 = ~(sub_487_2_n_10 | ~sub_487_2_n_79);
 assign sub_487_2_n_87 = ~sub_487_2_n_86;
 assign sub_487_2_n_85 = ~(sub_487_2_n_76 | ~sub_487_2_n_74);
 assign sub_487_2_n_84 = ~(sub_487_2_n_52 & (sub_487_2_n_44 | sub_487_2_n_3));
 assign sub_487_2_n_83 = ~(sub_487_2_n_55 & (sub_487_2_n_47 | sub_487_2_n_54));
 assign sub_487_2_n_88 = ~(sub_487_2_n_60 | sub_487_2_n_13);
 assign sub_487_2_n_86 = ~(sub_487_2_n_57 & (sub_487_2_n_38 | sub_487_2_n_2));
 assign sub_487_2_n_82 = ~sub_487_2_n_10;
 assign sub_487_2_n_80 = ~sub_487_2_n_79;
 assign sub_487_2_n_78 = ~sub_487_2_n_77;
 assign sub_487_2_n_76 = ~sub_487_2_n_75;
 assign sub_487_2_n_74 = ~(sub_487_2_n_54 & sub_487_2_n_55);
 assign sub_487_2_n_73 = ~(sub_487_2_n_49 | sub_487_2_n_56);
 assign sub_487_2_n_72 = (sub_487_2_n_50 | {in2[15]});
 assign sub_487_2_n_71 = ~(sub_487_2_n_3 | ~sub_487_2_n_52);
 assign sub_487_2_n_81 = ~(sub_487_2_n_13 | sub_487_2_n_48);
 assign sub_487_2_n_70 = ~(sub_487_2_n_49 & ~sub_487_2_n_8);
 assign sub_487_2_n_79 = ~(sub_487_2_n_1 | sub_487_2_n_2);
 assign sub_487_2_n_77 = ~(sub_487_2_n_8 | sub_487_2_n_56);
 assign sub_487_2_n_75 = ~(sub_487_2_n_5 | sub_487_2_n_48);
 assign sub_487_2_n_65 = ~sub_487_2_n_64;
 assign sub_487_2_n_63 = ~(sub_487_2_n_9 & ~sub_487_2_n_46);
 assign sub_487_2_n_62 = ~(sub_487_2_n_7 | sub_487_2_n_46);
 assign sub_487_2_n_61 = ~({in2[20]} | ({in2[21]} | ({in2[22]} | {in2[23]})));
 assign sub_487_2_n_60 = ~(sub_487_2_n_43 | sub_487_2_n_48);
 assign in1_43_0_ = ~(sub_487_2_n_53 & ~(sub_487_2_n_40 & {in1[34]}));
 assign sub_487_2_n_58 = ~({in2[16]} | ({in2[17]} | ({in2[18]} | {in2[19]})));
 assign sub_487_2_n_69 = ~(sub_487_2_n_6 | sub_487_2_n_3);
 assign sub_487_2_n_68 = ~(sub_487_2_n_12 | sub_487_2_n_56);
 assign sub_487_2_n_67 = ~(sub_487_2_n_14 | sub_487_2_n_54);
 assign sub_487_2_n_66 = ~(sub_487_2_n_45 & ~sub_487_2_n_7);
 assign sub_487_2_n_64 = ~(sub_487_2_n_11 | sub_487_2_n_0);
 assign sub_487_2_n_55 = ~sub_487_2_n_14;
 assign sub_487_2_n_54 = ~sub_487_2_n_9;
 assign sub_487_2_n_57 = ~(in1_41_12_ & ~{in2[13]});
 assign sub_487_2_n_38 = ~(in1_41_11_ & ~{in2[12]});
 assign sub_487_2_n_56 = ~(in1_41_6_ | sub_487_2_n_42);
 assign sub_487_2_n_53 = ~({in2[0]} & ~{in1[34]});
 assign sub_487_2_n_52 = ~(in1_41_10_ & ~{in2[11]});
 assign sub_487_2_n_51 = ~(in1_41_4_ & ~{in2[5]});
 assign sub_487_2_n_50 = ~(in1_41_13_ & ~{in2[14]});
 assign sub_487_2_n_37 = ~(in1_41_3_ & ~{in2[4]});
 assign sub_487_2_n_49 = ~(in1_41_5_ & ~{in2[6]});
 assign sub_487_2_n_48 = ~(in1_41_8_ | sub_487_2_n_41);
 assign sub_487_2_n_47 = ~(in1_41_1_ & ~{in2[2]});
 assign sub_487_2_n_46 = ~(in1_41_1_ | ~{in2[2]});
 assign sub_487_2_n_45 = ~(in1_41_0_ & ~{in2[1]});
 assign sub_487_2_n_44 = ~(in1_41_9_ & ~{in2[10]});
 assign sub_487_2_n_43 = ~(in1_41_7_ & ~{in2[8]});
 assign sub_487_2_n_42 = ~{in2[7]};
 assign sub_487_2_n_41 = ~{in2[9]};
 assign sub_487_2_n_40 = ~{in2[0]};
 assign in1_43_4_ = ~(sub_487_2_n_109 ^ sub_487_2_n_19);
 assign sub_487_2_n_35 = ~(sub_487_2_n_76 | ~sub_487_2_n_102);
 assign sub_487_2_n_34 = ~(sub_487_2_n_119 | ~sub_487_2_n_101);
 assign in1_43_10_ = ~(sub_487_2_n_118 ^ sub_487_2_n_16);
 assign in1_43_9_ = (sub_487_2_n_122 ^ sub_487_2_n_81);
 assign in1_43_8_ = ~(sub_487_2_n_117 ^ sub_487_2_n_15);
 assign in1_43_12_ = ~(sub_487_2_n_34 ^ sub_487_2_n_23);
 assign sub_487_2_n_29 = ~(sub_487_2_n_88 | ~sub_487_2_n_69);
 assign in1_43_7_ = (sub_487_2_n_121 ^ sub_487_2_n_68);
 assign in1_43_3_ = (sub_487_2_n_107 ^ sub_487_2_n_67);
 assign in1_43_5_ = (sub_487_2_n_114 ^ sub_487_2_n_21);
 assign in1_43_2_ = ~(sub_487_2_n_17 ^ sub_487_2_n_18);
 assign sub_487_2_n_24 = ~(sub_487_2_n_2 | ~sub_487_2_n_57);
 assign sub_487_2_n_23 = ~(sub_487_2_n_1 | ~sub_487_2_n_38);
 assign sub_487_2_n_22 = (sub_487_2_n_0 | (sub_487_2_n_37 & sub_487_2_n_51));
 assign sub_487_2_n_21 = ~(sub_487_2_n_0 | ~sub_487_2_n_51);
 assign sub_487_2_n_20 = (sub_487_2_n_50 & sub_487_2_n_4);
 assign sub_487_2_n_19 = ~(sub_487_2_n_11 | ~sub_487_2_n_37);
 assign sub_487_2_n_18 = ~(sub_487_2_n_46 | ~sub_487_2_n_47);
 assign sub_487_2_n_17 = ~(sub_487_2_n_100 | ~sub_487_2_n_45);
 assign sub_487_2_n_16 = ~(sub_487_2_n_6 | ~sub_487_2_n_44);
 assign sub_487_2_n_15 = ~(sub_487_2_n_5 | ~sub_487_2_n_43);
 assign sub_487_2_n_14 = ~({in2[3]} | ~in1_41_2_);
 assign sub_487_2_n_13 = (in1_41_8_ & sub_487_2_n_41);
 assign sub_487_2_n_12 = (in1_41_6_ & sub_487_2_n_42);
 assign sub_487_2_n_11 = ~(in1_41_3_ | ~{in2[4]});
 assign sub_487_2_n_10 = ~(sub_487_2_n_4 & ~{in2[15]});
 assign sub_487_2_n_9 = ~({in2[3]} & ~in1_41_2_);
 assign sub_487_2_n_8 = ~(in1_41_5_ | ~{in2[6]});
 assign sub_487_2_n_7 = ~(in1_41_0_ | ~{in2[1]});
 assign sub_487_2_n_6 = ~(in1_41_9_ | ~{in2[10]});
 assign sub_487_2_n_5 = ~(in1_41_7_ | ~{in2[8]});
 assign sub_487_2_n_4 = ~({in2[14]} & ~in1_41_13_);
 assign sub_487_2_n_3 = ~(in1_41_10_ | ~{in2[11]});
 assign sub_487_2_n_2 = ~(in1_41_12_ | ~{in2[13]});
 assign sub_487_2_n_1 = ~(in1_41_11_ | ~{in2[12]});
 assign sub_487_2_n_0 = ~(in1_41_4_ | ~{in2[5]});
 assign in1_46_15_ = ~(sub_508_2_n_154 & ~sub_508_2_n_155);
 assign sub_508_2_n_155 = ~(sub_508_2_n_42 | (sub_508_2_n_52 | sub_508_2_n_26));
 assign sub_508_2_n_154 = ~(sub_508_2_n_26 & (sub_508_2_n_42 | sub_508_2_n_52));
 assign in1_46_14_ = ~(sub_508_2_n_151 & ~sub_508_2_n_150);
 assign in1_46_13_ = ~(sub_508_2_n_149 & ~sub_508_2_n_148);
 assign sub_508_2_n_151 = ~(sub_508_2_n_146 & ~sub_508_2_n_94);
 assign sub_508_2_n_150 = ~(sub_508_2_n_146 | ~sub_508_2_n_94);
 assign sub_508_2_n_149 = ~(sub_508_2_n_41 & ~sub_508_2_n_28);
 assign sub_508_2_n_148 = ~(sub_508_2_n_143 | (sub_508_2_n_61 | ~sub_508_2_n_28));
 assign in1_46_24_ = ~(sub_508_2_n_140 & sub_508_2_n_103);
 assign sub_508_2_n_146 = ~(sub_508_2_n_108 & (sub_508_2_n_38 | sub_508_2_n_25));
 assign in1_46_9_ = ~(sub_508_2_n_141 & ~sub_508_2_n_142);
 assign in1_46_7_ = ~((sub_508_2_n_88 & ~sub_508_2_n_137) | (sub_508_2_n_22 & sub_508_2_n_137));
 assign sub_508_2_n_143 = ~(sub_508_2_n_38 | sub_508_2_n_58);
 assign sub_508_2_n_142 = ~(sub_508_2_n_138 | sub_508_2_n_20);
 assign sub_508_2_n_141 = ~(sub_508_2_n_138 & sub_508_2_n_20);
 assign sub_508_2_n_140 = ~(sub_508_2_n_37 & sub_508_2_n_127);
 assign sub_508_2_n_139 = ~(sub_508_2_n_71 & (sub_508_2_n_133 | sub_508_2_n_14));
 assign sub_508_2_n_138 = ~(sub_508_2_n_70 & (sub_508_2_n_131 | sub_508_2_n_11));
 assign sub_508_2_n_137 = ~(sub_508_2_n_68 | (sub_508_2_n_132 & sub_508_2_n_66));
 assign in1_46_10_ = ~(sub_508_2_n_133 ^ sub_508_2_n_27);
 assign in1_46_5_ = ~((sub_508_2_n_74 & ~sub_508_2_n_39) | (sub_508_2_n_75 & sub_508_2_n_39));
 assign sub_508_2_n_134 = ~(sub_508_2_n_131 | sub_508_2_n_102);
 assign sub_508_2_n_133 = ~(sub_508_2_n_123 | sub_508_2_n_130);
 assign sub_508_2_n_132 = ~(sub_508_2_n_43 & (sub_508_2_n_44 | sub_508_2_n_77));
 assign sub_508_2_n_131 = ~(sub_508_2_n_129 | sub_508_2_n_122);
 assign sub_508_2_n_130 = ~(sub_508_2_n_117 | sub_508_2_n_128);
 assign sub_508_2_n_129 = ~(sub_508_2_n_128 | sub_508_2_n_113);
 assign sub_508_2_n_128 = ~(sub_508_2_n_126 | sub_508_2_n_3);
 assign sub_508_2_n_127 = ~(sub_508_2_n_125 | sub_508_2_n_118);
 assign sub_508_2_n_44 = ~(sub_508_2_n_124 | sub_508_2_n_98);
 assign sub_508_2_n_126 = ~(sub_508_2_n_120 & sub_508_2_n_53);
 assign sub_508_2_n_125 = ~(sub_508_2_n_119 | sub_508_2_n_106);
 assign sub_508_2_n_124 = ~(sub_508_2_n_21 | sub_508_2_n_17);
 assign sub_508_2_n_123 = ~(sub_508_2_n_36 & sub_508_2_n_35);
 assign sub_508_2_n_122 = ~(sub_508_2_n_101 & (sub_508_2_n_43 | sub_508_2_n_91));
 assign in1_46_1_ = ~(sub_508_2_n_112 & ~sub_508_2_n_111);
 assign sub_508_2_n_120 = ~(sub_508_2_n_109 & sub_508_2_n_83);
 assign sub_508_2_n_119 = ~(sub_508_2_n_114 | sub_508_2_n_99);
 assign sub_508_2_n_118 = ~(sub_508_2_n_110 & sub_508_2_n_18);
 assign sub_508_2_n_117 = ~(sub_508_2_n_105 & sub_508_2_n_104);
 assign sub_508_2_n_116 = ~(sub_508_2_n_101 | sub_508_2_n_93);
 assign sub_508_2_n_115 = ~(sub_508_2_n_0 | ~sub_508_2_n_50);
 assign sub_508_2_n_114 = ~(sub_508_2_n_100 | sub_508_2_n_23);
 assign sub_508_2_n_113 = ~(sub_508_2_n_104 & sub_508_2_n_90);
 assign sub_508_2_n_112 = ~(sub_508_2_n_95 & sub_508_2_n_50);
 assign sub_508_2_n_111 = ~(sub_508_2_n_95 | sub_508_2_n_50);
 assign sub_508_2_n_110 = ~(sub_508_2_n_107 & sub_508_2_n_86);
 assign sub_508_2_n_109 = ~(sub_508_2_n_65 & ~sub_508_2_n_50);
 assign sub_508_2_n_108 = ~sub_508_2_n_107;
 assign sub_508_2_n_103 = (sub_508_2_n_79 & sub_508_2_n_80);
 assign sub_508_2_n_102 = ~(sub_508_2_n_92 & sub_508_2_n_76);
 assign sub_508_2_n_107 = ~(sub_508_2_n_73 & (sub_508_2_n_60 | sub_508_2_n_2));
 assign sub_508_2_n_106 = ~(sub_508_2_n_86 & ~sub_508_2_n_25);
 assign sub_508_2_n_105 = ~(sub_508_2_n_91 | sub_508_2_n_93);
 assign sub_508_2_n_104 = (sub_508_2_n_78 & sub_508_2_n_1);
 assign sub_508_2_n_99 = ~(sub_508_2_n_63 & (sub_508_2_n_71 | sub_508_2_n_12));
 assign sub_508_2_n_98 = ~(sub_508_2_n_72 & (sub_508_2_n_53 | sub_508_2_n_64));
 assign sub_508_2_n_101 = ~(sub_508_2_n_89 | sub_508_2_n_6);
 assign sub_508_2_n_100 = ~(sub_508_2_n_82 | sub_508_2_n_5);
 assign sub_508_2_n_43 = ~(sub_508_2_n_84 | sub_508_2_n_13);
 assign sub_508_2_n_93 = ~sub_508_2_n_92;
 assign sub_508_2_n_91 = ~sub_508_2_n_90;
 assign sub_508_2_n_89 = ~(sub_508_2_n_67 | sub_508_2_n_69);
 assign sub_508_2_n_97 = ~(sub_508_2_n_61 | sub_508_2_n_58);
 assign sub_508_2_n_96 = ~(sub_508_2_n_3 | sub_508_2_n_64);
 assign sub_508_2_n_95 = ~(sub_508_2_n_65 & ~sub_508_2_n_0);
 assign sub_508_2_n_88 = ~(sub_508_2_n_6 | sub_508_2_n_69);
 assign sub_508_2_n_94 = ~(sub_508_2_n_52 | sub_508_2_n_15);
 assign sub_508_2_n_92 = ~(sub_508_2_n_11 | sub_508_2_n_59);
 assign sub_508_2_n_90 = ~(sub_508_2_n_8 | sub_508_2_n_69);
 assign sub_508_2_n_84 = ~(sub_508_2_n_56 | sub_508_2_n_55);
 assign sub_508_2_n_83 = ~(sub_508_2_n_0 | sub_508_2_n_9);
 assign sub_508_2_n_82 = ~(sub_508_2_n_70 | sub_508_2_n_59);
 assign in1_46_0_ = ~(sub_508_2_n_50 & ~(sub_508_2_n_47 & {in1[33]}));
 assign sub_508_2_n_80 = ~({in2[20]} | ({in2[21]} | ({in2[22]} | {in2[23]})));
 assign sub_508_2_n_79 = ~({in2[16]} | ({in2[17]} | ({in2[18]} | {in2[19]})));
 assign sub_508_2_n_87 = ~(sub_508_2_n_68 | sub_508_2_n_8);
 assign sub_508_2_n_86 = ~(sub_508_2_n_15 | sub_508_2_n_7);
 assign sub_508_2_n_78 = ~(sub_508_2_n_4 | sub_508_2_n_55);
 assign sub_508_2_n_77 = ~(sub_508_2_n_54 & ~sub_508_2_n_4);
 assign sub_508_2_n_85 = ~(sub_508_2_n_57 | sub_508_2_n_4);
 assign sub_508_2_n_76 = ~(sub_508_2_n_14 | sub_508_2_n_12);
 assign sub_508_2_n_75 = ~(sub_508_2_n_54 & ~sub_508_2_n_13);
 assign sub_508_2_n_74 = ~(sub_508_2_n_13 | sub_508_2_n_55);
 assign sub_508_2_n_72 = ~sub_508_2_n_3;
 assign sub_508_2_n_68 = ~sub_508_2_n_67;
 assign sub_508_2_n_66 = ~sub_508_2_n_8;
 assign sub_508_2_n_64 = ~sub_508_2_n_1;
 assign sub_508_2_n_73 = ~(in1_44_12_ & ~{in2[13]});
 assign sub_508_2_n_71 = ~(in1_44_9_ & ~{in2[10]});
 assign sub_508_2_n_70 = ~(in1_44_7_ & ~{in2[8]});
 assign sub_508_2_n_69 = ~(in1_44_6_ | sub_508_2_n_48);
 assign sub_508_2_n_67 = ~(in1_44_5_ & ~{in2[6]});
 assign sub_508_2_n_65 = ~(in1_44_0_ & ~{in2[1]});
 assign sub_508_2_n_61 = ~sub_508_2_n_60;
 assign sub_508_2_n_58 = ~sub_508_2_n_10;
 assign sub_508_2_n_57 = ~sub_508_2_n_56;
 assign sub_508_2_n_54 = ~sub_508_2_n_55;
 assign sub_508_2_n_52 = ~sub_508_2_n_51;
 assign sub_508_2_n_63 = ~(in1_44_10_ & ~{in2[11]});
 assign sub_508_2_n_62 = ~(in1_44_14_ & ~{in2[15]});
 assign sub_508_2_n_60 = ~(in1_44_11_ & ~{in2[12]});
 assign sub_508_2_n_59 = ~(in1_44_8_ | sub_508_2_n_46);
 assign sub_508_2_n_56 = ~(in1_44_3_ & ~{in2[4]});
 assign sub_508_2_n_55 = ~(in1_44_4_ | sub_508_2_n_49);
 assign sub_508_2_n_53 = ~(in1_44_1_ & ~{in2[2]});
 assign sub_508_2_n_51 = ~(in1_44_13_ & ~{in2[14]});
 assign sub_508_2_n_50 = ~({in2[0]} & ~{in1[33]});
 assign sub_508_2_n_49 = ~{in2[5]};
 assign sub_508_2_n_48 = ~{in2[7]};
 assign sub_508_2_n_47 = ~{in2[0]};
 assign sub_508_2_n_46 = ~{in2[9]};
 assign sub_508_2_n_42 = ~(sub_508_2_n_15 | ~sub_508_2_n_146);
 assign sub_508_2_n_41 = (sub_508_2_n_143 | sub_508_2_n_61);
 assign in1_46_6_ = (sub_508_2_n_132 ^ sub_508_2_n_87);
 assign sub_508_2_n_39 = ~(sub_508_2_n_57 | ~(sub_508_2_n_44 | sub_508_2_n_4));
 assign sub_508_2_n_38 = ~(sub_508_2_n_134 | ~sub_508_2_n_119);
 assign sub_508_2_n_37 = ~(sub_508_2_n_134 & ~sub_508_2_n_106);
 assign sub_508_2_n_36 = ~(sub_508_2_n_116 | ~sub_508_2_n_100);
 assign sub_508_2_n_35 = ~(sub_508_2_n_105 & ~sub_508_2_n_43);
 assign in1_46_12_ = ~(sub_508_2_n_38 ^ sub_508_2_n_97);
 assign in1_46_3_ = (sub_508_2_n_126 ^ sub_508_2_n_96);
 assign in1_46_11_ = (sub_508_2_n_139 ^ sub_508_2_n_19);
 assign in1_46_2_ = ~(sub_508_2_n_21 ^ sub_508_2_n_16);
 assign in1_46_8_ = ~(sub_508_2_n_131 ^ sub_508_2_n_24);
 assign in1_46_4_ = ~(sub_508_2_n_44 ^ sub_508_2_n_85);
 assign sub_508_2_n_28 = ~(sub_508_2_n_2 | ~sub_508_2_n_73);
 assign sub_508_2_n_27 = ~(sub_508_2_n_14 | ~sub_508_2_n_71);
 assign sub_508_2_n_26 = ~(sub_508_2_n_62 & ~sub_508_2_n_7);
 assign sub_508_2_n_25 = ~(sub_508_2_n_10 & ~sub_508_2_n_2);
 assign sub_508_2_n_24 = ~(sub_508_2_n_11 | ~sub_508_2_n_70);
 assign sub_508_2_n_23 = (sub_508_2_n_12 | sub_508_2_n_14);
 assign sub_508_2_n_22 = (sub_508_2_n_69 | sub_508_2_n_6);
 assign sub_508_2_n_21 = ~(sub_508_2_n_115 | ~sub_508_2_n_65);
 assign sub_508_2_n_20 = (sub_508_2_n_5 | sub_508_2_n_59);
 assign sub_508_2_n_19 = ~(sub_508_2_n_12 | ~sub_508_2_n_63);
 assign sub_508_2_n_18 = (sub_508_2_n_62 & (sub_508_2_n_51 | sub_508_2_n_7));
 assign sub_508_2_n_17 = ~(sub_508_2_n_1 & ~sub_508_2_n_9);
 assign sub_508_2_n_16 = ~(sub_508_2_n_9 | ~sub_508_2_n_53);
 assign sub_508_2_n_15 = ~(in1_44_13_ | ~{in2[14]});
 assign sub_508_2_n_14 = ~(in1_44_9_ | ~{in2[10]});
 assign sub_508_2_n_13 = (in1_44_4_ & sub_508_2_n_49);
 assign sub_508_2_n_12 = ~(in1_44_10_ | ~{in2[11]});
 assign sub_508_2_n_11 = ~(in1_44_7_ | ~{in2[8]});
 assign sub_508_2_n_10 = ~({in2[12]} & ~in1_44_11_);
 assign sub_508_2_n_9 = ~(in1_44_1_ | ~{in2[2]});
 assign sub_508_2_n_8 = ~(in1_44_5_ | ~{in2[6]});
 assign sub_508_2_n_7 = ~(in1_44_14_ | ~{in2[15]});
 assign sub_508_2_n_6 = (in1_44_6_ & sub_508_2_n_48);
 assign sub_508_2_n_5 = (in1_44_8_ & sub_508_2_n_46);
 assign sub_508_2_n_4 = ~(in1_44_3_ | ~{in2[4]});
 assign sub_508_2_n_3 = ~({in2[3]} | ~in1_44_2_);
 assign sub_508_2_n_2 = ~(in1_44_12_ | ~{in2[13]});
 assign sub_508_2_n_1 = ~({in2[3]} & ~in1_44_2_);
 assign sub_508_2_n_0 = ~(in1_44_0_ | ~{in2[1]});
 assign in1_49_11_ = ~(sub_529_2_n_154 & ~sub_529_2_n_155);
 assign sub_529_2_n_155 = ~(sub_529_2_n_152 | sub_529_2_n_27);
 assign sub_529_2_n_154 = ~(sub_529_2_n_152 & sub_529_2_n_27);
 assign sub_529_2_n_153 = ~(sub_529_2_n_48 & (sub_529_2_n_151 | sub_529_2_n_4));
 assign sub_529_2_n_152 = ~(sub_529_2_n_65 | (sub_529_2_n_145 & sub_529_2_n_71));
 assign sub_529_2_n_151 = ~sub_529_2_n_150;
 assign sub_529_2_n_150 = ~(sub_529_2_n_102 & (sub_529_2_n_140 | sub_529_2_n_23));
 assign sub_529_2_n_149 = ~(sub_529_2_n_58 & (sub_529_2_n_140 | sub_529_2_n_70));
 assign in1_49_24_ = ~sub_529_2_n_147;
 assign sub_529_2_n_147 = ~(sub_529_2_n_146 | sub_529_2_n_133);
 assign sub_529_2_n_146 = ~(sub_529_2_n_141 | sub_529_2_n_132);
 assign sub_529_2_n_145 = ~(sub_529_2_n_105 & (sub_529_2_n_136 | sub_529_2_n_89));
 assign sub_529_2_n_144 = ~(sub_529_2_n_50 & (sub_529_2_n_136 | sub_529_2_n_6));
 assign sub_529_2_n_143 = ~(sub_529_2_n_51 & (sub_529_2_n_139 | sub_529_2_n_46));
 assign sub_529_2_n_142 = ~(sub_529_2_n_43 & (sub_529_2_n_136 | sub_529_2_n_116));
 assign sub_529_2_n_141 = ~(sub_529_2_n_136 | sub_529_2_n_99);
 assign sub_529_2_n_140 = ~(sub_529_2_n_134 | (sub_529_2_n_124 | sub_529_2_n_117));
 assign sub_529_2_n_139 = ~sub_529_2_n_138;
 assign sub_529_2_n_138 = ~(sub_529_2_n_98 & (sub_529_2_n_130 | sub_529_2_n_19));
 assign sub_529_2_n_137 = ~(sub_529_2_n_69 & (sub_529_2_n_130 | sub_529_2_n_68));
 assign sub_529_2_n_136 = ~(sub_529_2_n_135 | sub_529_2_n_122);
 assign sub_529_2_n_135 = ~(sub_529_2_n_111 | sub_529_2_n_13);
 assign sub_529_2_n_134 = ~(sub_529_2_n_41 | sub_529_2_n_13);
 assign sub_529_2_n_133 = ~(sub_529_2_n_115 & (sub_529_2_n_121 | sub_529_2_n_110));
 assign sub_529_2_n_132 = ~(sub_529_2_n_125 & sub_529_2_n_120);
 assign in1_49_2_ = ~(sub_529_2_n_127 & ~sub_529_2_n_128);
 assign sub_529_2_n_130 = ~(sub_529_2_n_126 | sub_529_2_n_95);
 assign sub_529_2_n_129 = ~(sub_529_2_n_118 & sub_529_2_n_59);
 assign sub_529_2_n_128 = ~(sub_529_2_n_119 | sub_529_2_n_17);
 assign sub_529_2_n_127 = ~(sub_529_2_n_119 & sub_529_2_n_17);
 assign sub_529_2_n_126 = ~(sub_529_2_n_119 | sub_529_2_n_18);
 assign sub_529_2_n_125 = ~(sub_529_2_n_117 | sub_529_2_n_114);
 assign sub_529_2_n_124 = ~(sub_529_2_n_123 & sub_529_2_n_112);
 assign sub_529_2_n_123 = ~(sub_529_2_n_106 & sub_529_2_n_100);
 assign sub_529_2_n_122 = ~(sub_529_2_n_103 & (sub_529_2_n_98 | sub_529_2_n_16));
 assign sub_529_2_n_121 = ~(sub_529_2_n_85 | (sub_529_2_n_102 & sub_529_2_n_23));
 assign sub_529_2_n_120 = (sub_529_2_n_109 & sub_529_2_n_96);
 assign sub_529_2_n_119 = ~(sub_529_2_n_113 | sub_529_2_n_61);
 assign sub_529_2_n_118 = ~(sub_529_2_n_108 & sub_529_2_n_83);
 assign sub_529_2_n_117 = ~(sub_529_2_n_107 & sub_529_2_n_94);
 assign sub_529_2_n_116 = ~(sub_529_2_n_33 & ~sub_529_2_n_99);
 assign sub_529_2_n_115 = ~(sub_529_2_n_10 | ~sub_529_2_n_97);
 assign sub_529_2_n_114 = ~(sub_529_2_n_63 | ~sub_529_2_n_97);
 assign sub_529_2_n_113 = ~(sub_529_2_n_0 | ~sub_529_2_n_57);
 assign sub_529_2_n_112 = ~(sub_529_2_n_100 & ~sub_529_2_n_103);
 assign sub_529_2_n_110 = ~(sub_529_2_n_96 & sub_529_2_n_63);
 assign sub_529_2_n_109 = ~(sub_529_2_n_101 & sub_529_2_n_84);
 assign sub_529_2_n_108 = ~(sub_529_2_n_60 & ~sub_529_2_n_57);
 assign sub_529_2_n_107 = ~(sub_529_2_n_104 & sub_529_2_n_92);
 assign sub_529_2_n_111 = ~(sub_529_2_n_93 & sub_529_2_n_75);
 assign sub_529_2_n_106 = ~(sub_529_2_n_98 | sub_529_2_n_16);
 assign sub_529_2_n_105 = ~sub_529_2_n_104;
 assign sub_529_2_n_102 = ~sub_529_2_n_101;
 assign sub_529_2_n_99 = ~sub_529_2_n_100;
 assign sub_529_2_n_104 = ~(sub_529_2_n_73 & (sub_529_2_n_50 | sub_529_2_n_11));
 assign sub_529_2_n_103 = ~(sub_529_2_n_1 | ~(sub_529_2_n_51 | sub_529_2_n_49));
 assign sub_529_2_n_101 = ~(sub_529_2_n_67 & (sub_529_2_n_58 | sub_529_2_n_12));
 assign sub_529_2_n_100 = (sub_529_2_n_88 & sub_529_2_n_92);
 assign sub_529_2_n_95 = ~(sub_529_2_n_47 & (sub_529_2_n_59 | sub_529_2_n_9));
 assign sub_529_2_n_94 = ~(sub_529_2_n_78 | sub_529_2_n_74);
 assign sub_529_2_n_93 = (sub_529_2_n_79 & sub_529_2_n_76);
 assign sub_529_2_n_98 = ~(sub_529_2_n_8 | ~(sub_529_2_n_69 | sub_529_2_n_62));
 assign sub_529_2_n_97 = ~({in2[18]} | ({in2[19]} | ({in2[23]} | sub_529_2_n_81)));
 assign sub_529_2_n_96 = ~(sub_529_2_n_7 | ~(sub_529_2_n_48 | sub_529_2_n_72));
 assign sub_529_2_n_89 = ~sub_529_2_n_88;
 assign sub_529_2_n_85 = ~sub_529_2_n_84;
 assign sub_529_2_n_83 = ~(sub_529_2_n_0 | sub_529_2_n_5);
 assign sub_529_2_n_92 = ~(sub_529_2_n_3 | sub_529_2_n_66);
 assign sub_529_2_n_91 = ~(sub_529_2_n_1 | sub_529_2_n_49);
 assign sub_529_2_n_90 = ~(sub_529_2_n_7 | sub_529_2_n_72);
 assign sub_529_2_n_88 = ~(sub_529_2_n_6 | sub_529_2_n_11);
 assign sub_529_2_n_87 = ~(sub_529_2_n_65 | sub_529_2_n_3);
 assign sub_529_2_n_86 = ~(sub_529_2_n_47 & ~sub_529_2_n_9);
 assign sub_529_2_n_84 = ~(sub_529_2_n_4 | sub_529_2_n_72);
 assign sub_529_2_n_81 = ({in2[17]} | ({in2[20]} | ({in2[21]} | {in2[22]})));
 assign in1_49_0_ = ~(sub_529_2_n_57 & ~(sub_529_2_n_53 & {in1[32]}));
 assign sub_529_2_n_79 = ~(sub_529_2_n_9 & sub_529_2_n_47);
 assign sub_529_2_n_78 = ~(sub_529_2_n_64 | sub_529_2_n_66);
 assign sub_529_2_n_77 = ~(sub_529_2_n_61 | sub_529_2_n_0);
 assign sub_529_2_n_76 = ~(sub_529_2_n_68 | sub_529_2_n_62);
 assign sub_529_2_n_75 = ~(sub_529_2_n_46 | sub_529_2_n_49);
 assign sub_529_2_n_82 = ~(sub_529_2_n_8 | sub_529_2_n_62);
 assign sub_529_2_n_71 = ~sub_529_2_n_3;
 assign sub_529_2_n_70 = ~sub_529_2_n_2;
 assign sub_529_2_n_74 = (sub_529_2_n_55 & in1_47_10_);
 assign sub_529_2_n_73 = ~(in1_47_8_ & ~{in2[9]});
 assign sub_529_2_n_72 = ~(in1_47_14_ | ~{in2[15]});
 assign sub_529_2_n_51 = ~(in1_47_5_ & ~{in2[6]});
 assign sub_529_2_n_50 = ~(in1_47_7_ & ~{in2[8]});
 assign sub_529_2_n_69 = ~(in1_47_3_ & ~{in2[4]});
 assign sub_529_2_n_68 = ~(in1_47_3_ | ~{in2[4]});
 assign sub_529_2_n_65 = ~sub_529_2_n_64;
 assign sub_529_2_n_61 = ~sub_529_2_n_60;
 assign sub_529_2_n_67 = ~(in1_47_12_ & ~{in2[13]});
 assign sub_529_2_n_66 = ~(in1_47_10_ | sub_529_2_n_55);
 assign sub_529_2_n_64 = ~(in1_47_9_ & ~{in2[10]});
 assign sub_529_2_n_63 = ~(in1_47_15_ & ~{in2[16]});
 assign sub_529_2_n_62 = ~(in1_47_4_ | ~{in2[5]});
 assign sub_529_2_n_60 = ~(in1_47_0_ & ~{in2[1]});
 assign sub_529_2_n_59 = ~(in1_47_1_ & ~{in2[2]});
 assign sub_529_2_n_49 = ~(in1_47_6_ | sub_529_2_n_54);
 assign sub_529_2_n_48 = ~(in1_47_13_ & ~{in2[14]});
 assign sub_529_2_n_58 = ~(in1_47_11_ & ~{in2[12]});
 assign sub_529_2_n_47 = ~(in1_47_2_ & ~{in2[3]});
 assign sub_529_2_n_57 = ~({in2[0]} & ~{in1[32]});
 assign sub_529_2_n_56 = ~{in2[6]};
 assign sub_529_2_n_55 = ~{in2[11]};
 assign sub_529_2_n_54 = ~{in2[7]};
 assign sub_529_2_n_53 = ~{in2[0]};
 assign sub_529_2_n_46 = ~(in1_47_5_ | sub_529_2_n_56);
 assign in1_49_10_ = (sub_529_2_n_145 ^ sub_529_2_n_87);
 assign in1_49_3_ = ~(sub_529_2_n_129 ^ sub_529_2_n_86);
 assign sub_529_2_n_43 = ~(sub_529_2_n_42 | ~sub_529_2_n_120);
 assign sub_529_2_n_42 = (sub_529_2_n_117 & sub_529_2_n_33);
 assign sub_529_2_n_41 = ~(sub_529_2_n_100 & ~sub_529_2_n_111);
 assign in1_49_1_ = (sub_529_2_n_77 ^ sub_529_2_n_57);
 assign in1_49_13_ = (sub_529_2_n_149 ^ sub_529_2_n_21);
 assign in1_49_16_ = (sub_529_2_n_142 ^ sub_529_2_n_20);
 assign in1_49_7_ = (sub_529_2_n_143 ^ sub_529_2_n_91);
 assign in1_49_15_ = (sub_529_2_n_153 ^ sub_529_2_n_90);
 assign in1_49_14_ = (sub_529_2_n_150 ^ sub_529_2_n_15);
 assign in1_49_12_ = ~(sub_529_2_n_140 ^ sub_529_2_n_14);
 assign sub_529_2_n_33 = ~(sub_529_2_n_85 | sub_529_2_n_23);
 assign in1_49_8_ = ~(sub_529_2_n_136 ^ sub_529_2_n_24);
 assign in1_49_6_ = (sub_529_2_n_138 ^ sub_529_2_n_25);
 assign in1_49_4_ = ~(sub_529_2_n_130 ^ sub_529_2_n_22);
 assign in1_49_5_ = (sub_529_2_n_137 ^ sub_529_2_n_82);
 assign in1_49_9_ = (sub_529_2_n_144 ^ sub_529_2_n_26);
 assign sub_529_2_n_27 = ~(sub_529_2_n_66 | sub_529_2_n_74);
 assign sub_529_2_n_26 = ~(sub_529_2_n_11 | ~sub_529_2_n_73);
 assign sub_529_2_n_25 = ~(sub_529_2_n_46 | ~sub_529_2_n_51);
 assign sub_529_2_n_24 = ~(sub_529_2_n_6 | ~sub_529_2_n_50);
 assign sub_529_2_n_23 = ~(sub_529_2_n_2 & ~sub_529_2_n_12);
 assign sub_529_2_n_22 = ~(sub_529_2_n_68 | ~sub_529_2_n_69);
 assign sub_529_2_n_21 = ~(sub_529_2_n_12 | ~sub_529_2_n_67);
 assign sub_529_2_n_20 = ~(sub_529_2_n_10 | ~sub_529_2_n_63);
 assign sub_529_2_n_19 = (sub_529_2_n_62 | sub_529_2_n_68);
 assign sub_529_2_n_18 = (sub_529_2_n_5 | sub_529_2_n_9);
 assign sub_529_2_n_17 = ~(sub_529_2_n_5 | ~sub_529_2_n_59);
 assign sub_529_2_n_16 = (sub_529_2_n_49 | sub_529_2_n_46);
 assign sub_529_2_n_15 = ~(sub_529_2_n_4 | ~sub_529_2_n_48);
 assign sub_529_2_n_14 = ~(sub_529_2_n_70 | ~sub_529_2_n_58);
 assign sub_529_2_n_13 = ~(sub_529_2_n_129 | ~sub_529_2_n_47);
 assign sub_529_2_n_12 = ~(in1_47_12_ | ~{in2[13]});
 assign sub_529_2_n_11 = ~(in1_47_8_ | ~{in2[9]});
 assign sub_529_2_n_10 = ~(in1_47_15_ | ~{in2[16]});
 assign sub_529_2_n_9 = ~(in1_47_2_ | ~{in2[3]});
 assign sub_529_2_n_8 = ~({in2[5]} | ~in1_47_4_);
 assign sub_529_2_n_7 = ~({in2[15]} | ~in1_47_14_);
 assign sub_529_2_n_6 = ~(in1_47_7_ | ~{in2[8]});
 assign sub_529_2_n_5 = ~(in1_47_1_ | ~{in2[2]});
 assign sub_529_2_n_4 = ~(in1_47_13_ | ~{in2[14]});
 assign sub_529_2_n_3 = ~(in1_47_9_ | ~{in2[10]});
 assign sub_529_2_n_2 = ~({in2[12]} & ~in1_47_11_);
 assign sub_529_2_n_1 = (in1_47_6_ & sub_529_2_n_54);
 assign sub_529_2_n_0 = ~(in1_47_0_ | ~{in2[1]});
 assign in1_52_15_ = (sub_550_2_n_148 ^ sub_550_2_n_28);
 assign in1_52_17_ = (sub_550_2_n_144 ^ sub_550_2_n_89);
 assign sub_550_2_n_148 = ~(sub_550_2_n_65 & (sub_550_2_n_142 | sub_550_2_n_0));
 assign in1_52_14_ = (sub_550_2_n_141 ^ sub_550_2_n_23);
 assign in1_52_13_ = (sub_550_2_n_140 ^ sub_550_2_n_86);
 assign in1_52_24_ = (sub_550_2_n_138 & sub_550_2_n_111);
 assign sub_550_2_n_144 = ~(sub_550_2_n_70 & (sub_550_2_n_136 | sub_550_2_n_69));
 assign in1_52_16_ = ~(sub_550_2_n_136 ^ sub_550_2_n_26);
 assign sub_550_2_n_142 = ~sub_550_2_n_141;
 assign sub_550_2_n_141 = ~(sub_550_2_n_101 & (sub_550_2_n_135 | sub_550_2_n_95));
 assign sub_550_2_n_140 = ~(sub_550_2_n_61 & (sub_550_2_n_135 | sub_550_2_n_12));
 assign sub_550_2_n_139 = ~(sub_550_2_n_62 & (sub_550_2_n_38 | sub_550_2_n_10));
 assign sub_550_2_n_138 = ~(sub_550_2_n_117 & (sub_550_2_n_134 | sub_550_2_n_114));
 assign in1_52_9_ = (sub_550_2_n_133 ^ sub_550_2_n_74);
 assign sub_550_2_n_136 = ~(sub_550_2_n_118 | (sub_550_2_n_131 & sub_550_2_n_104));
 assign sub_550_2_n_135 = ~sub_550_2_n_134;
 assign sub_550_2_n_134 = ~(sub_550_2_n_112 & (sub_550_2_n_130 | sub_550_2_n_107));
 assign sub_550_2_n_133 = ~(sub_550_2_n_57 & (sub_550_2_n_130 | sub_550_2_n_11));
 assign sub_550_2_n_132 = ~(sub_550_2_n_59 & (sub_550_2_n_129 | sub_550_2_n_6));
 assign sub_550_2_n_131 = ~(sub_550_2_n_130 | sub_550_2_n_107);
 assign sub_550_2_n_130 = ~(sub_550_2_n_126 | sub_550_2_n_113);
 assign sub_550_2_n_129 = ~sub_550_2_n_128;
 assign sub_550_2_n_128 = ~(sub_550_2_n_100 & (sub_550_2_n_124 | sub_550_2_n_24));
 assign sub_550_2_n_127 = ~(sub_550_2_n_60 & (sub_550_2_n_124 | sub_550_2_n_15));
 assign sub_550_2_n_126 = ~(sub_550_2_n_108 | sub_550_2_n_125);
 assign sub_550_2_n_125 = ~(sub_550_2_n_122 | sub_550_2_n_44);
 assign sub_550_2_n_124 = ~(sub_550_2_n_123 | sub_550_2_n_99);
 assign sub_550_2_n_123 = ~(sub_550_2_n_41 | sub_550_2_n_3);
 assign sub_550_2_n_122 = ~(sub_550_2_n_58 & (sub_550_2_n_46 | sub_550_2_n_1));
 assign in1_52_2_ = ~(sub_550_2_n_119 & ~sub_550_2_n_120);
 assign sub_550_2_n_120 = ~(sub_550_2_n_46 | sub_550_2_n_18);
 assign sub_550_2_n_119 = ~(sub_550_2_n_46 & sub_550_2_n_18);
 assign sub_550_2_n_118 = ~(sub_550_2_n_116 & sub_550_2_n_45);
 assign sub_550_2_n_117 = ~(sub_550_2_n_115 | (sub_550_2_n_45 & sub_550_2_n_103));
 assign sub_550_2_n_116 = ~(sub_550_2_n_104 & ~sub_550_2_n_112);
 assign sub_550_2_n_115 = ~(sub_550_2_n_7 & ~sub_550_2_n_39);
 assign sub_550_2_n_114 = ~sub_550_2_n_45;
 assign sub_550_2_n_45 = ~(sub_550_2_n_109 | sub_550_2_n_98);
 assign sub_550_2_n_113 = ~(sub_550_2_n_97 & (sub_550_2_n_100 | sub_550_2_n_83));
 assign sub_550_2_n_112 = ~(sub_550_2_n_110 | sub_550_2_n_96);
 assign sub_550_2_n_46 = ~(sub_550_2_n_40 | sub_550_2_n_67);
 assign sub_550_2_n_111 = ~(sub_550_2_n_106 & (sub_550_2_n_79 | sub_550_2_n_72));
 assign sub_550_2_n_110 = ~(sub_550_2_n_105 | sub_550_2_n_25);
 assign sub_550_2_n_109 = ~(sub_550_2_n_101 | sub_550_2_n_16);
 assign sub_550_2_n_108 = ~(sub_550_2_n_102 & sub_550_2_n_78);
 assign sub_550_2_n_104 = ~sub_550_2_n_103;
 assign sub_550_2_n_107 = ~(sub_550_2_n_84 & sub_550_2_n_88);
 assign sub_550_2_n_102 = (sub_550_2_n_87 & sub_550_2_n_82);
 assign sub_550_2_n_106 = ~({in2[22]} | ({in2[23]} | ~sub_550_2_n_76));
 assign sub_550_2_n_105 = ~(sub_550_2_n_90 | sub_550_2_n_14);
 assign sub_550_2_n_103 = ~(sub_550_2_n_94 & sub_550_2_n_75);
 assign sub_550_2_n_99 = ~(sub_550_2_n_43 & (sub_550_2_n_58 | sub_550_2_n_3));
 assign sub_550_2_n_98 = ~(sub_550_2_n_73 & (sub_550_2_n_65 | sub_550_2_n_8));
 assign sub_550_2_n_97 = ~(sub_550_2_n_81 | sub_550_2_n_9);
 assign sub_550_2_n_96 = ~(sub_550_2_n_71 & (sub_550_2_n_62 | sub_550_2_n_13));
 assign sub_550_2_n_101 = ~(sub_550_2_n_80 | sub_550_2_n_5);
 assign sub_550_2_n_100 = ~(sub_550_2_n_91 | sub_550_2_n_4);
 assign sub_550_2_n_95 = ~sub_550_2_n_94;
 assign sub_550_2_n_91 = ~(sub_550_2_n_60 | sub_550_2_n_66);
 assign sub_550_2_n_90 = ~(sub_550_2_n_57 | sub_550_2_n_63);
 assign sub_550_2_n_89 = ~(sub_550_2_n_72 | sub_550_2_n_56);
 assign sub_550_2_n_94 = ~(sub_550_2_n_12 | sub_550_2_n_68);
 assign sub_550_2_n_93 = ~(sub_550_2_n_44 | sub_550_2_n_3);
 assign sub_550_2_n_88 = ~(sub_550_2_n_10 | sub_550_2_n_13);
 assign sub_550_2_n_92 = ~(sub_550_2_n_4 | sub_550_2_n_66);
 assign sub_550_2_n_87 = ~(sub_550_2_n_15 | sub_550_2_n_66);
 assign sub_550_2_n_86 = ~(sub_550_2_n_5 | sub_550_2_n_68);
 assign sub_550_2_n_83 = ~sub_550_2_n_82;
 assign sub_550_2_n_81 = ~(sub_550_2_n_59 | sub_550_2_n_64);
 assign sub_550_2_n_80 = ~(sub_550_2_n_61 | sub_550_2_n_68);
 assign sub_550_2_n_79 = ~(sub_550_2_n_70 | sub_550_2_n_56);
 assign sub_550_2_n_78 = ~(sub_550_2_n_3 & sub_550_2_n_43);
 assign in1_52_0_ = ~(sub_550_2_n_54 & ~(sub_550_2_n_49 & {in1[31]}));
 assign sub_550_2_n_76 = ~({in2[18]} | ({in2[19]} | ({in2[20]} | {in2[21]})));
 assign sub_550_2_n_85 = ~(sub_550_2_n_9 | sub_550_2_n_64);
 assign sub_550_2_n_84 = ~(sub_550_2_n_11 | sub_550_2_n_63);
 assign sub_550_2_n_75 = ~(sub_550_2_n_0 | sub_550_2_n_8);
 assign sub_550_2_n_74 = ~(sub_550_2_n_14 | sub_550_2_n_63);
 assign sub_550_2_n_82 = ~(sub_550_2_n_6 | sub_550_2_n_64);
 assign sub_550_2_n_69 = ~sub_550_2_n_7;
 assign sub_550_2_n_44 = ~sub_550_2_n_43;
 assign sub_550_2_n_73 = ~(in1_50_14_ & ~{in2[15]});
 assign sub_550_2_n_72 = (sub_550_2_n_51 & in1_50_16_);
 assign sub_550_2_n_71 = ~(in1_50_10_ & ~{in2[11]});
 assign sub_550_2_n_67 = ~(sub_550_2_n_48 | ~sub_550_2_n_53);
 assign sub_550_2_n_70 = ~(in1_50_15_ & ~{in2[16]});
 assign sub_550_2_n_68 = ~(in1_50_12_ | ~{in2[13]});
 assign sub_550_2_n_43 = ~(in1_50_2_ & ~{in2[3]});
 assign sub_550_2_n_56 = ~sub_550_2_n_55;
 assign sub_550_2_n_66 = ~(in1_50_4_ | ~{in2[5]});
 assign sub_550_2_n_65 = ~(in1_50_13_ & ~{in2[14]});
 assign sub_550_2_n_64 = ~(in1_50_6_ | sub_550_2_n_50);
 assign sub_550_2_n_63 = ~(in1_50_8_ | sub_550_2_n_52);
 assign sub_550_2_n_62 = ~(in1_50_9_ & ~{in2[10]});
 assign sub_550_2_n_61 = ~(in1_50_11_ & ~{in2[12]});
 assign sub_550_2_n_60 = ~(in1_50_3_ & ~{in2[4]});
 assign sub_550_2_n_59 = ~(in1_50_5_ & ~{in2[6]});
 assign sub_550_2_n_58 = ~(in1_50_1_ & ~{in2[2]});
 assign sub_550_2_n_57 = ~(in1_50_7_ & ~{in2[8]});
 assign sub_550_2_n_55 = (in1_50_16_ | sub_550_2_n_51);
 assign sub_550_2_n_54 = ~({in2[0]} & ~{in1[31]});
 assign sub_550_2_n_53 = ~{in2[1]};
 assign sub_550_2_n_52 = ~{in2[9]};
 assign sub_550_2_n_51 = ~{in2[17]};
 assign sub_550_2_n_50 = ~{in2[7]};
 assign sub_550_2_n_49 = ~{in2[0]};
 assign sub_550_2_n_48 = ~in1_50_0_;
 assign in1_52_10_ = ~(sub_550_2_n_38 ^ sub_550_2_n_22);
 assign sub_550_2_n_41 = (sub_550_2_n_46 | sub_550_2_n_1);
 assign sub_550_2_n_40 = (sub_550_2_n_54 & (in1_50_0_ | sub_550_2_n_53));
 assign sub_550_2_n_39 = ~(sub_550_2_n_55 & sub_550_2_n_106);
 assign sub_550_2_n_38 = ~(sub_550_2_n_30 | ~sub_550_2_n_105);
 assign in1_52_8_ = ~(sub_550_2_n_130 ^ sub_550_2_n_17);
 assign in1_52_3_ = (sub_550_2_n_122 ^ sub_550_2_n_93);
 assign in1_52_5_ = (sub_550_2_n_127 ^ sub_550_2_n_92);
 assign in1_52_12_ = ~(sub_550_2_n_135 ^ sub_550_2_n_21);
 assign in1_52_11_ = (sub_550_2_n_139 ^ sub_550_2_n_27);
 assign in1_52_4_ = ~(sub_550_2_n_124 ^ sub_550_2_n_20);
 assign in1_52_7_ = (sub_550_2_n_132 ^ sub_550_2_n_85);
 assign sub_550_2_n_30 = ~(sub_550_2_n_130 | ~sub_550_2_n_84);
 assign in1_52_6_ = (sub_550_2_n_128 ^ sub_550_2_n_19);
 assign sub_550_2_n_28 = ~(sub_550_2_n_8 | ~sub_550_2_n_73);
 assign sub_550_2_n_27 = ~(sub_550_2_n_13 | ~sub_550_2_n_71);
 assign sub_550_2_n_26 = ~(sub_550_2_n_69 | ~sub_550_2_n_70);
 assign sub_550_2_n_25 = (sub_550_2_n_13 | sub_550_2_n_10);
 assign sub_550_2_n_24 = (sub_550_2_n_66 | sub_550_2_n_15);
 assign sub_550_2_n_23 = ~(sub_550_2_n_0 | ~sub_550_2_n_65);
 assign sub_550_2_n_22 = ~(sub_550_2_n_10 | ~sub_550_2_n_62);
 assign sub_550_2_n_21 = ~(sub_550_2_n_12 | ~sub_550_2_n_61);
 assign sub_550_2_n_20 = ~(sub_550_2_n_15 | ~sub_550_2_n_60);
 assign sub_550_2_n_19 = ~(sub_550_2_n_6 | ~sub_550_2_n_59);
 assign sub_550_2_n_18 = ~(sub_550_2_n_1 | ~sub_550_2_n_58);
 assign sub_550_2_n_17 = ~(sub_550_2_n_11 | ~sub_550_2_n_57);
 assign sub_550_2_n_16 = (sub_550_2_n_8 | sub_550_2_n_0);
 assign sub_550_2_n_15 = ~(in1_50_3_ | ~{in2[4]});
 assign sub_550_2_n_14 = (in1_50_8_ & sub_550_2_n_52);
 assign sub_550_2_n_13 = ~(in1_50_10_ | ~{in2[11]});
 assign sub_550_2_n_12 = ~(in1_50_11_ | ~{in2[12]});
 assign sub_550_2_n_11 = ~(in1_50_7_ | ~{in2[8]});
 assign sub_550_2_n_10 = ~(in1_50_9_ | ~{in2[10]});
 assign sub_550_2_n_9 = (in1_50_6_ & sub_550_2_n_50);
 assign sub_550_2_n_8 = ~(in1_50_14_ | ~{in2[15]});
 assign sub_550_2_n_7 = ~({in2[16]} & ~in1_50_15_);
 assign sub_550_2_n_6 = ~(in1_50_5_ | ~{in2[6]});
 assign sub_550_2_n_5 = ~({in2[13]} | ~in1_50_12_);
 assign sub_550_2_n_4 = ~({in2[5]} | ~in1_50_4_);
 assign sub_550_2_n_3 = ~(in1_50_2_ | ~{in2[3]});
 assign sub_550_2_n_1 = ~(in1_50_1_ | ~{in2[2]});
 assign sub_550_2_n_0 = ~(in1_50_13_ | ~{in2[14]});
 assign in1_52_1_ = (sub_550_2_n_48 ^ ({in2[1]} ^ sub_550_2_n_54));
 assign in1_55_18_ = ~(sub_571_2_n_143 ^ sub_571_2_n_20);
 assign sub_571_2_n_146 = ~(sub_571_2_n_69 & (sub_571_2_n_139 | sub_571_2_n_11));
 assign in1_55_24_ = ~(sub_571_2_n_142 | sub_571_2_n_122);
 assign in1_55_14_ = ~((sub_571_2_n_18 & ~sub_571_2_n_139) | (sub_571_2_n_101 & sub_571_2_n_139));
 assign sub_571_2_n_143 = ~(sub_571_2_n_115 & (sub_571_2_n_136 | sub_571_2_n_17));
 assign sub_571_2_n_142 = ~(sub_571_2_n_136 | (sub_571_2_n_17 | sub_571_2_n_113));
 assign sub_571_2_n_141 = ~(sub_571_2_n_79 & (sub_571_2_n_136 | sub_571_2_n_62));
 assign in1_55_16_ = ~(sub_571_2_n_136 ^ sub_571_2_n_26);
 assign sub_571_2_n_139 = ~(sub_571_2_n_110 | (sub_571_2_n_134 & sub_571_2_n_95));
 assign sub_571_2_n_138 = ~(sub_571_2_n_73 & (sub_571_2_n_48 | sub_571_2_n_9));
 assign sub_571_2_n_137 = ~(sub_571_2_n_78 & (sub_571_2_n_46 | sub_571_2_n_5));
 assign sub_571_2_n_136 = ~(sub_571_2_n_135 | sub_571_2_n_123);
 assign sub_571_2_n_135 = ~(sub_571_2_n_130 | (sub_571_2_n_116 | sub_571_2_n_114));
 assign sub_571_2_n_134 = ~sub_571_2_n_48;
 assign sub_571_2_n_133 = ~(sub_571_2_n_75 & (sub_571_2_n_130 | sub_571_2_n_64));
 assign sub_571_2_n_132 = ~(sub_571_2_n_130 | sub_571_2_n_116);
 assign sub_571_2_n_131 = ~(sub_571_2_n_81 | (sub_571_2_n_128 & sub_571_2_n_67));
 assign sub_571_2_n_130 = ~(sub_571_2_n_129 | sub_571_2_n_119);
 assign sub_571_2_n_129 = ~(sub_571_2_n_125 | (sub_571_2_n_19 | sub_571_2_n_23));
 assign sub_571_2_n_128 = ~(sub_571_2_n_111 & (sub_571_2_n_125 | sub_571_2_n_19));
 assign sub_571_2_n_127 = ~(sub_571_2_n_65 & (sub_571_2_n_125 | sub_571_2_n_77));
 assign sub_571_2_n_126 = ~(sub_571_2_n_52 & (sub_571_2_n_117 | sub_571_2_n_68));
 assign sub_571_2_n_125 = ~(sub_571_2_n_124 | sub_571_2_n_106);
 assign sub_571_2_n_124 = ~(sub_571_2_n_117 | sub_571_2_n_15);
 assign sub_571_2_n_123 = ~(sub_571_2_n_120 & (sub_571_2_n_118 | sub_571_2_n_114));
 assign sub_571_2_n_122 = ~(sub_571_2_n_121 | sub_571_2_n_91);
 assign sub_571_2_n_121 = ~(sub_571_2_n_43 | sub_571_2_n_97);
 assign sub_571_2_n_120 = ~(sub_571_2_n_30 | sub_571_2_n_112);
 assign sub_571_2_n_119 = ~(sub_571_2_n_107 & (sub_571_2_n_111 | sub_571_2_n_23));
 assign sub_571_2_n_118 = ~(sub_571_2_n_44 | sub_571_2_n_105);
 assign sub_571_2_n_117 = ~(sub_571_2_n_47 | sub_571_2_n_72);
 assign sub_571_2_n_116 = ~(sub_571_2_n_99 & sub_571_2_n_104);
 assign sub_571_2_n_113 = ~(sub_571_2_n_103 & ~sub_571_2_n_91);
 assign sub_571_2_n_112 = ~(sub_571_2_n_70 & (sub_571_2_n_69 | sub_571_2_n_13));
 assign sub_571_2_n_115 = ~(sub_571_2_n_89 | ~sub_571_2_n_83);
 assign sub_571_2_n_114 = ~(sub_571_2_n_95 & sub_571_2_n_90);
 assign sub_571_2_n_110 = ~sub_571_2_n_109;
 assign sub_571_2_n_107 = ~(sub_571_2_n_87 | sub_571_2_n_4);
 assign sub_571_2_n_106 = ~(sub_571_2_n_82 & (sub_571_2_n_52 | sub_571_2_n_12));
 assign sub_571_2_n_105 = ~(sub_571_2_n_84 & (sub_571_2_n_78 | sub_571_2_n_8));
 assign sub_571_2_n_111 = ~(sub_571_2_n_86 | sub_571_2_n_6);
 assign sub_571_2_n_109 = ~(sub_571_2_n_96 | sub_571_2_n_2);
 assign sub_571_2_n_108 = ~(sub_571_2_n_98 | sub_571_2_n_3);
 assign sub_571_2_n_101 = ~sub_571_2_n_18;
 assign sub_571_2_n_98 = ~(sub_571_2_n_75 | sub_571_2_n_76);
 assign sub_571_2_n_97 = ~(sub_571_2_n_71 | {in2[19]});
 assign sub_571_2_n_96 = ~(sub_571_2_n_73 | sub_571_2_n_63);
 assign sub_571_2_n_104 = ~(sub_571_2_n_5 | sub_571_2_n_8);
 assign sub_571_2_n_103 = ~(sub_571_2_n_14 | {in2[19]});
 assign sub_571_2_n_102 = ~(sub_571_2_n_6 | sub_571_2_n_51);
 assign sub_571_2_n_100 = ~(sub_571_2_n_2 | sub_571_2_n_63);
 assign sub_571_2_n_99 = ~(sub_571_2_n_64 | sub_571_2_n_76);
 assign sub_571_2_n_89 = ~(sub_571_2_n_79 | sub_571_2_n_0);
 assign in1_55_0_ = ~(sub_571_2_n_61 & ~(sub_571_2_n_54 & {in1[30]}));
 assign sub_571_2_n_87 = ~(sub_571_2_n_80 | sub_571_2_n_74);
 assign sub_571_2_n_86 = ~(sub_571_2_n_65 | sub_571_2_n_51);
 assign sub_571_2_n_95 = ~(sub_571_2_n_9 | sub_571_2_n_63);
 assign sub_571_2_n_94 = ~(sub_571_2_n_4 | sub_571_2_n_74);
 assign sub_571_2_n_85 = ~(sub_571_2_n_78 & ~sub_571_2_n_5);
 assign sub_571_2_n_93 = ~(sub_571_2_n_3 | sub_571_2_n_76);
 assign sub_571_2_n_92 = ~(sub_571_2_n_81 | sub_571_2_n_66);
 assign sub_571_2_n_91 = ({in2[20]} | ({in2[21]} | ({in2[22]} | {in2[23]})));
 assign sub_571_2_n_90 = ~(sub_571_2_n_11 | sub_571_2_n_13);
 assign sub_571_2_n_81 = ~sub_571_2_n_80;
 assign sub_571_2_n_77 = ~sub_571_2_n_10;
 assign sub_571_2_n_84 = ~(in1_53_10_ & ~{in2[11]});
 assign sub_571_2_n_83 = ~(in1_53_16_ & ~{in2[17]});
 assign sub_571_2_n_82 = ~(in1_53_2_ & ~{in2[3]});
 assign sub_571_2_n_72 = ~(sub_571_2_n_57 | ~sub_571_2_n_56);
 assign sub_571_2_n_80 = ~(in1_53_5_ & ~{in2[6]});
 assign sub_571_2_n_79 = ~(in1_53_15_ & ~{in2[16]});
 assign sub_571_2_n_78 = ~(in1_53_9_ & ~{in2[10]});
 assign sub_571_2_n_52 = ~(in1_53_1_ & ~{in2[2]});
 assign sub_571_2_n_76 = ~(in1_53_8_ | sub_571_2_n_55);
 assign sub_571_2_n_75 = ~(in1_53_7_ & ~{in2[8]});
 assign sub_571_2_n_74 = ~(in1_53_6_ | sub_571_2_n_58);
 assign sub_571_2_n_73 = ~(in1_53_11_ & ~{in2[12]});
 assign sub_571_2_n_67 = ~sub_571_2_n_66;
 assign sub_571_2_n_62 = ~sub_571_2_n_1;
 assign sub_571_2_n_71 = ~(in1_53_17_ & ~{in2[18]});
 assign sub_571_2_n_70 = ~(in1_53_14_ & ~{in2[15]});
 assign sub_571_2_n_51 = ~(in1_53_4_ | sub_571_2_n_60);
 assign sub_571_2_n_69 = ~(in1_53_13_ & ~{in2[14]});
 assign sub_571_2_n_68 = ~(in1_53_1_ | ~{in2[2]});
 assign sub_571_2_n_66 = ~(in1_53_5_ | ~{in2[6]});
 assign sub_571_2_n_65 = ~(in1_53_3_ & ~{in2[4]});
 assign sub_571_2_n_64 = ~(in1_53_7_ | ~{in2[8]});
 assign sub_571_2_n_63 = ~(in1_53_12_ | sub_571_2_n_59);
 assign sub_571_2_n_61 = ~({in2[0]} & ~{in1[30]});
 assign sub_571_2_n_60 = ~{in2[5]};
 assign sub_571_2_n_59 = ~{in2[13]};
 assign sub_571_2_n_58 = ~{in2[7]};
 assign sub_571_2_n_57 = ~in1_53_0_;
 assign sub_571_2_n_56 = ~{in2[1]};
 assign sub_571_2_n_55 = ~{in2[9]};
 assign sub_571_2_n_54 = ~{in2[0]};
 assign in1_55_10_ = (sub_571_2_n_46 ^ sub_571_2_n_85);
 assign in1_55_6_ = (sub_571_2_n_128 ^ sub_571_2_n_92);
 assign sub_571_2_n_48 = ~(sub_571_2_n_132 | ~sub_571_2_n_118);
 assign sub_571_2_n_47 = (sub_571_2_n_61 & (in1_53_0_ | sub_571_2_n_56));
 assign sub_571_2_n_46 = ~(sub_571_2_n_38 | ~sub_571_2_n_108);
 assign in1_55_17_ = (sub_571_2_n_141 ^ sub_571_2_n_28);
 assign sub_571_2_n_44 = ~(sub_571_2_n_108 | ~sub_571_2_n_104);
 assign sub_571_2_n_43 = ~(sub_571_2_n_115 | ~sub_571_2_n_103);
 assign in1_55_15_ = (sub_571_2_n_146 ^ sub_571_2_n_21);
 assign in1_55_5_ = (sub_571_2_n_127 ^ sub_571_2_n_102);
 assign in1_55_13_ = (sub_571_2_n_138 ^ sub_571_2_n_100);
 assign in1_55_2_ = ~(sub_571_2_n_117 ^ sub_571_2_n_25);
 assign sub_571_2_n_38 = ~(sub_571_2_n_130 | ~sub_571_2_n_99);
 assign in1_55_12_ = ~(sub_571_2_n_48 ^ sub_571_2_n_22);
 assign in1_55_11_ = (sub_571_2_n_137 ^ sub_571_2_n_29);
 assign in1_55_7_ = ~(sub_571_2_n_131 ^ sub_571_2_n_94);
 assign in1_55_8_ = ~(sub_571_2_n_130 ^ sub_571_2_n_24);
 assign in1_55_4_ = ~(sub_571_2_n_125 ^ sub_571_2_n_16);
 assign in1_55_3_ = (sub_571_2_n_126 ^ sub_571_2_n_27);
 assign in1_55_9_ = (sub_571_2_n_133 ^ sub_571_2_n_93);
 assign sub_571_2_n_30 = ~(sub_571_2_n_109 | ~sub_571_2_n_90);
 assign sub_571_2_n_29 = ~(sub_571_2_n_8 | ~sub_571_2_n_84);
 assign sub_571_2_n_28 = ~(sub_571_2_n_0 | ~sub_571_2_n_83);
 assign sub_571_2_n_27 = ~(sub_571_2_n_12 | ~sub_571_2_n_82);
 assign sub_571_2_n_26 = ~(sub_571_2_n_62 | ~sub_571_2_n_79);
 assign sub_571_2_n_25 = ~(sub_571_2_n_68 | ~sub_571_2_n_52);
 assign sub_571_2_n_24 = ~(sub_571_2_n_64 | ~sub_571_2_n_75);
 assign sub_571_2_n_23 = (sub_571_2_n_74 | sub_571_2_n_66);
 assign sub_571_2_n_22 = ~(sub_571_2_n_9 | ~sub_571_2_n_73);
 assign sub_571_2_n_21 = ~(sub_571_2_n_13 | ~sub_571_2_n_70);
 assign sub_571_2_n_20 = ~(sub_571_2_n_71 & ~sub_571_2_n_14);
 assign sub_571_2_n_19 = ~(sub_571_2_n_10 & ~sub_571_2_n_51);
 assign sub_571_2_n_18 = ~(sub_571_2_n_11 | ~sub_571_2_n_69);
 assign sub_571_2_n_17 = ~(sub_571_2_n_1 & ~sub_571_2_n_0);
 assign sub_571_2_n_16 = ~(sub_571_2_n_77 | ~sub_571_2_n_65);
 assign sub_571_2_n_15 = (sub_571_2_n_12 | sub_571_2_n_68);
 assign sub_571_2_n_14 = ~(in1_53_17_ | ~{in2[18]});
 assign sub_571_2_n_13 = ~(in1_53_14_ | ~{in2[15]});
 assign sub_571_2_n_12 = ~(in1_53_2_ | ~{in2[3]});
 assign sub_571_2_n_11 = ~(in1_53_13_ | ~{in2[14]});
 assign sub_571_2_n_10 = ~({in2[4]} & ~in1_53_3_);
 assign sub_571_2_n_9 = ~(in1_53_11_ | ~{in2[12]});
 assign sub_571_2_n_8 = ~(in1_53_10_ | ~{in2[11]});
 assign sub_571_2_n_6 = (in1_53_4_ & sub_571_2_n_60);
 assign sub_571_2_n_5 = ~(in1_53_9_ | ~{in2[10]});
 assign sub_571_2_n_4 = (in1_53_6_ & sub_571_2_n_58);
 assign sub_571_2_n_3 = (in1_53_8_ & sub_571_2_n_55);
 assign sub_571_2_n_2 = (in1_53_12_ & sub_571_2_n_59);
 assign sub_571_2_n_1 = ~({in2[16]} & ~in1_53_15_);
 assign sub_571_2_n_0 = ~(in1_53_16_ | ~{in2[17]});
 assign in1_55_1_ = (sub_571_2_n_57 ^ ({in2[1]} ^ sub_571_2_n_61));
 assign in1_58_19_ = ~(sub_592_2_n_162 ^ sub_592_2_n_24);
 assign sub_592_2_n_162 = ~(sub_592_2_n_161 | sub_592_2_n_81);
 assign sub_592_2_n_161 = ~(sub_592_2_n_46 | sub_592_2_n_0);
 assign in1_58_13_ = (sub_592_2_n_154 ^ sub_592_2_n_17);
 assign in1_58_24_ = ~(sub_592_2_n_158 | sub_592_2_n_137);
 assign sub_592_2_n_158 = ~(sub_592_2_n_156 | sub_592_2_n_38);
 assign sub_592_2_n_157 = ~(sub_592_2_n_84 & (sub_592_2_n_152 | sub_592_2_n_12));
 assign sub_592_2_n_156 = ~(sub_592_2_n_151 & sub_592_2_n_104);
 assign sub_592_2_n_155 = ~(sub_592_2_n_120 | ~(sub_592_2_n_150 | sub_592_2_n_99));
 assign sub_592_2_n_154 = ~(sub_592_2_n_79 | ~(sub_592_2_n_150 | sub_592_2_n_8));
 assign sub_592_2_n_153 = ~(sub_592_2_n_67 & (sub_592_2_n_43 | sub_592_2_n_48));
 assign sub_592_2_n_152 = ~sub_592_2_n_151;
 assign sub_592_2_n_151 = ~(sub_592_2_n_138 & (sub_592_2_n_146 | (sub_592_2_n_31 | sub_592_2_n_123)));
 assign sub_592_2_n_150 = ~(sub_592_2_n_135 | (sub_592_2_n_145 & sub_592_2_n_125));
 assign sub_592_2_n_149 = ~(sub_592_2_n_68 & (sub_592_2_n_146 | sub_592_2_n_1));
 assign in1_58_8_ = ~(sub_592_2_n_145 ^ sub_592_2_n_89);
 assign sub_592_2_n_147 = ~(sub_592_2_n_83 & (sub_592_2_n_143 | sub_592_2_n_72));
 assign sub_592_2_n_145 = ~sub_592_2_n_146;
 assign sub_592_2_n_146 = ~(sub_592_2_n_144 | sub_592_2_n_131);
 assign sub_592_2_n_144 = ~(sub_592_2_n_51 | (sub_592_2_n_15 | sub_592_2_n_19));
 assign sub_592_2_n_143 = ~(sub_592_2_n_118 | (sub_592_2_n_140 & sub_592_2_n_112));
 assign sub_592_2_n_142 = ~(sub_592_2_n_64 | (sub_592_2_n_140 & sub_592_2_n_3));
 assign sub_592_2_n_141 = ~(sub_592_2_n_85 & (sub_592_2_n_130 | sub_592_2_n_82));
 assign sub_592_2_n_140 = ~sub_592_2_n_51;
 assign sub_592_2_n_51 = ~(sub_592_2_n_139 | sub_592_2_n_113);
 assign sub_592_2_n_139 = ~(sub_592_2_n_130 | sub_592_2_n_13);
 assign sub_592_2_n_138 = ~(sub_592_2_n_136 | sub_592_2_n_133);
 assign sub_592_2_n_137 = ~(sub_592_2_n_132 | sub_592_2_n_95);
 assign sub_592_2_n_136 = ~(sub_592_2_n_134 | sub_592_2_n_123);
 assign sub_592_2_n_135 = ~sub_592_2_n_134;
 assign sub_592_2_n_134 = ~(sub_592_2_n_127 | sub_592_2_n_121);
 assign sub_592_2_n_133 = ~(sub_592_2_n_122 & (sub_592_2_n_119 | sub_592_2_n_97));
 assign sub_592_2_n_132 = ~(sub_592_2_n_126 | sub_592_2_n_115);
 assign sub_592_2_n_131 = ~(sub_592_2_n_114 & (sub_592_2_n_117 | sub_592_2_n_19));
 assign sub_592_2_n_130 = ~(sub_592_2_n_128 | sub_592_2_n_4);
 assign in1_58_1_ = ~(in1_56_0_ ^ ({in2[1]} ^ sub_592_2_n_77));
 assign sub_592_2_n_128 = ~(sub_592_2_n_76 | ~sub_592_2_n_77);
 assign sub_592_2_n_127 = ~(sub_592_2_n_124 | sub_592_2_n_14);
 assign sub_592_2_n_126 = ~(sub_592_2_n_116 | sub_592_2_n_23);
 assign sub_592_2_n_125 = ~sub_592_2_n_31;
 assign sub_592_2_n_122 = ~(sub_592_2_n_105 | sub_592_2_n_10);
 assign sub_592_2_n_121 = ~(sub_592_2_n_88 & (sub_592_2_n_67 | sub_592_2_n_5));
 assign sub_592_2_n_124 = ~(sub_592_2_n_87 | ~(sub_592_2_n_68 | sub_592_2_n_47));
 assign sub_592_2_n_123 = ~(sub_592_2_n_98 & sub_592_2_n_96);
 assign sub_592_2_n_120 = ~sub_592_2_n_119;
 assign sub_592_2_n_118 = ~sub_592_2_n_117;
 assign sub_592_2_n_115 = ~(sub_592_2_n_86 & (sub_592_2_n_80 | sub_592_2_n_9));
 assign sub_592_2_n_114 = ~(sub_592_2_n_91 | sub_592_2_n_2);
 assign sub_592_2_n_113 = ~(sub_592_2_n_75 & (sub_592_2_n_85 | sub_592_2_n_11));
 assign sub_592_2_n_119 = ~(sub_592_2_n_92 | sub_592_2_n_74);
 assign sub_592_2_n_117 = ~(sub_592_2_n_90 | sub_592_2_n_6);
 assign sub_592_2_n_116 = ~(sub_592_2_n_94 | sub_592_2_n_73);
 assign sub_592_2_n_112 = ~sub_592_2_n_15;
 assign sub_592_2_n_105 = ~(sub_592_2_n_69 | ~sub_592_2_n_71);
 assign sub_592_2_n_104 = ~(sub_592_2_n_12 | sub_592_2_n_65);
 assign sub_592_2_n_111 = ~(sub_592_2_n_81 | sub_592_2_n_0);
 assign sub_592_2_n_110 = ~(sub_592_2_n_73 | sub_592_2_n_65);
 assign sub_592_2_n_109 = ~(sub_592_2_n_10 | sub_592_2_n_69);
 assign sub_592_2_n_108 = ~(sub_592_2_n_71 | sub_592_2_n_66);
 assign sub_592_2_n_107 = ~(sub_592_2_n_1 | sub_592_2_n_47);
 assign sub_592_2_n_106 = ~(sub_592_2_n_2 | sub_592_2_n_50);
 assign sub_592_2_n_99 = ~sub_592_2_n_98;
 assign sub_592_2_n_97 = ~sub_592_2_n_96;
 assign sub_592_2_n_94 = ~(sub_592_2_n_84 | sub_592_2_n_65);
 assign in1_58_0_ = ~(sub_592_2_n_77 & ~(sub_592_2_n_62 & {in1[29]}));
 assign sub_592_2_n_92 = ~(sub_592_2_n_78 | sub_592_2_n_70);
 assign sub_592_2_n_91 = ~(sub_592_2_n_50 | ~sub_592_2_n_7);
 assign sub_592_2_n_90 = ~(sub_592_2_n_63 | sub_592_2_n_49);
 assign sub_592_2_n_103 = ~(sub_592_2_n_6 | sub_592_2_n_49);
 assign sub_592_2_n_102 = ~(sub_592_2_n_87 | sub_592_2_n_47);
 assign sub_592_2_n_89 = ~(sub_592_2_n_68 & ~sub_592_2_n_1);
 assign sub_592_2_n_101 = ~(sub_592_2_n_79 | sub_592_2_n_8);
 assign sub_592_2_n_100 = ~(sub_592_2_n_7 | sub_592_2_n_72);
 assign sub_592_2_n_98 = ~(sub_592_2_n_8 | sub_592_2_n_70);
 assign sub_592_2_n_96 = ~(sub_592_2_n_66 | sub_592_2_n_69);
 assign sub_592_2_n_95 = ({in2[20]} | ({in2[21]} | ({in2[22]} | {in2[23]})));
 assign sub_592_2_n_83 = ~sub_592_2_n_7;
 assign sub_592_2_n_81 = ~sub_592_2_n_80;
 assign sub_592_2_n_79 = ~sub_592_2_n_78;
 assign sub_592_2_n_88 = ~(in1_56_10_ & ~{in2[11]});
 assign sub_592_2_n_76 = ~(in1_56_0_ | ~{in2[1]});
 assign sub_592_2_n_87 = (sub_592_2_n_53 & in1_56_8_);
 assign sub_592_2_n_86 = ~(in1_56_18_ & ~{in2[19]});
 assign sub_592_2_n_85 = ~(in1_56_1_ & ~{in2[2]});
 assign sub_592_2_n_84 = ~(in1_56_15_ & ~{in2[16]});
 assign sub_592_2_n_50 = ~(in1_56_6_ | sub_592_2_n_59);
 assign sub_592_2_n_82 = ~(in1_56_1_ | ~{in2[2]});
 assign sub_592_2_n_80 = ~(in1_56_17_ & ~{in2[18]});
 assign sub_592_2_n_78 = ~(in1_56_11_ & ~{in2[12]});
 assign sub_592_2_n_77 = ~({in2[0]} & ~{in1[29]});
 assign sub_592_2_n_64 = ~sub_592_2_n_63;
 assign sub_592_2_n_75 = ~(in1_56_2_ & ~{in2[3]});
 assign sub_592_2_n_74 = (sub_592_2_n_60 & in1_56_12_);
 assign sub_592_2_n_73 = (sub_592_2_n_55 & in1_56_16_);
 assign sub_592_2_n_72 = ~(in1_56_5_ | sub_592_2_n_56);
 assign sub_592_2_n_71 = (sub_592_2_n_58 & in1_56_13_);
 assign sub_592_2_n_70 = ~(in1_56_12_ | sub_592_2_n_60);
 assign sub_592_2_n_69 = ~(in1_56_14_ | sub_592_2_n_54);
 assign sub_592_2_n_68 = ~(in1_56_7_ & ~{in2[8]});
 assign sub_592_2_n_67 = ~(in1_56_9_ & ~{in2[10]});
 assign sub_592_2_n_66 = ~(in1_56_13_ | sub_592_2_n_58);
 assign sub_592_2_n_65 = ~(in1_56_16_ | sub_592_2_n_55);
 assign sub_592_2_n_49 = ~(in1_56_4_ | sub_592_2_n_57);
 assign sub_592_2_n_63 = ~(in1_56_3_ & ~{in2[4]});
 assign sub_592_2_n_62 = ~{in2[0]};
 assign sub_592_2_n_61 = ~{in2[10]};
 assign sub_592_2_n_60 = ~{in2[13]};
 assign sub_592_2_n_59 = ~{in2[7]};
 assign sub_592_2_n_58 = ~{in2[14]};
 assign sub_592_2_n_57 = ~{in2[5]};
 assign sub_592_2_n_56 = ~{in2[6]};
 assign sub_592_2_n_55 = ~{in2[17]};
 assign sub_592_2_n_54 = ~{in2[15]};
 assign sub_592_2_n_53 = ~{in2[9]};
 assign sub_592_2_n_48 = ~(in1_56_9_ | sub_592_2_n_61);
 assign sub_592_2_n_47 = ~(in1_56_8_ | sub_592_2_n_53);
 assign sub_592_2_n_46 = (sub_592_2_n_156 & sub_592_2_n_116);
 assign sub_592_2_n_45 = ~(sub_592_2_n_71 | ~(sub_592_2_n_155 | sub_592_2_n_66));
 assign in1_58_2_ = ~(sub_592_2_n_130 ^ sub_592_2_n_22);
 assign sub_592_2_n_43 = ~(sub_592_2_n_36 | ~sub_592_2_n_124);
 assign in1_58_18_ = ~(sub_592_2_n_46 ^ sub_592_2_n_111);
 assign in1_58_17_ = (sub_592_2_n_157 ^ sub_592_2_n_110);
 assign in1_58_16_ = (sub_592_2_n_151 ^ sub_592_2_n_20);
 assign in1_58_15_ = ~(sub_592_2_n_45 ^ sub_592_2_n_109);
 assign sub_592_2_n_38 = (sub_592_2_n_23 | sub_592_2_n_95);
 assign in1_58_14_ = ~(sub_592_2_n_155 ^ sub_592_2_n_108);
 assign sub_592_2_n_36 = ~(sub_592_2_n_146 | ~sub_592_2_n_107);
 assign in1_58_7_ = (sub_592_2_n_147 ^ sub_592_2_n_106);
 assign in1_58_4_ = ~(sub_592_2_n_51 ^ sub_592_2_n_21);
 assign in1_58_5_ = ~(sub_592_2_n_142 ^ sub_592_2_n_103);
 assign in1_58_9_ = (sub_592_2_n_149 ^ sub_592_2_n_102);
 assign sub_592_2_n_31 = ~(sub_592_2_n_107 & ~sub_592_2_n_14);
 assign in1_58_12_ = ~(sub_592_2_n_150 ^ sub_592_2_n_101);
 assign in1_58_6_ = ~(sub_592_2_n_143 ^ sub_592_2_n_100);
 assign in1_58_3_ = (sub_592_2_n_141 ^ sub_592_2_n_18);
 assign in1_58_10_ = ~(sub_592_2_n_43 ^ sub_592_2_n_16);
 assign in1_58_11_ = (sub_592_2_n_153 ^ sub_592_2_n_25);
 assign sub_592_2_n_25 = ~(sub_592_2_n_5 | ~sub_592_2_n_88);
 assign sub_592_2_n_24 = ~(sub_592_2_n_9 | ~sub_592_2_n_86);
 assign sub_592_2_n_23 = (sub_592_2_n_9 | sub_592_2_n_0);
 assign sub_592_2_n_22 = ~(sub_592_2_n_82 | ~sub_592_2_n_85);
 assign sub_592_2_n_21 = ~(sub_592_2_n_64 | ~sub_592_2_n_3);
 assign sub_592_2_n_20 = ~(sub_592_2_n_12 | ~sub_592_2_n_84);
 assign sub_592_2_n_19 = (sub_592_2_n_50 | sub_592_2_n_72);
 assign sub_592_2_n_18 = ~(sub_592_2_n_11 | ~sub_592_2_n_75);
 assign sub_592_2_n_17 = (sub_592_2_n_74 | sub_592_2_n_70);
 assign sub_592_2_n_16 = ~(sub_592_2_n_48 | ~sub_592_2_n_67);
 assign sub_592_2_n_15 = ~(sub_592_2_n_3 & ~sub_592_2_n_49);
 assign sub_592_2_n_14 = (sub_592_2_n_5 | sub_592_2_n_48);
 assign sub_592_2_n_13 = (sub_592_2_n_11 | sub_592_2_n_82);
 assign sub_592_2_n_12 = ~(in1_56_15_ | ~{in2[16]});
 assign sub_592_2_n_11 = ~(in1_56_2_ | ~{in2[3]});
 assign sub_592_2_n_10 = (in1_56_14_ & sub_592_2_n_54);
 assign sub_592_2_n_9 = ~(in1_56_18_ | ~{in2[19]});
 assign sub_592_2_n_8 = ~(in1_56_11_ | ~{in2[12]});
 assign sub_592_2_n_7 = (in1_56_5_ & sub_592_2_n_56);
 assign sub_592_2_n_6 = (in1_56_4_ & sub_592_2_n_57);
 assign sub_592_2_n_5 = ~(in1_56_10_ | ~{in2[11]});
 assign sub_592_2_n_4 = ~({in2[1]} | ~in1_56_0_);
 assign sub_592_2_n_3 = ~({in2[4]} & ~in1_56_3_);
 assign sub_592_2_n_2 = (in1_56_6_ & sub_592_2_n_59);
 assign sub_592_2_n_1 = ~(in1_56_7_ | ~{in2[8]});
 assign sub_592_2_n_0 = ~(in1_56_17_ | ~{in2[18]});
 assign in1_61_19_ = (sub_613_2_n_176 ^ sub_613_2_n_23);
 assign in1_61_15_ = ~((sub_613_2_n_114 & ~sub_613_2_n_44) | (sub_613_2_n_115 & sub_613_2_n_44));
 assign sub_613_2_n_176 = ~(sub_613_2_n_67 | ~(sub_613_2_n_173 | sub_613_2_n_13));
 assign in1_61_18_ = ~(sub_613_2_n_173 ^ sub_613_2_n_93);
 assign in1_61_24_ = ~(sub_613_2_n_172 | sub_613_2_n_149);
 assign sub_613_2_n_172 = ~(sub_613_2_n_167 | sub_613_2_n_132);
 assign sub_613_2_n_171 = ~(sub_613_2_n_86 | (sub_613_2_n_162 & sub_613_2_n_63));
 assign sub_613_2_n_173 = ~(sub_613_2_n_127 | (sub_613_2_n_162 & sub_613_2_n_116));
 assign in1_61_16_ = ~(sub_613_2_n_162 ^ sub_613_2_n_109);
 assign sub_613_2_n_169 = ~(sub_613_2_n_65 | (sub_613_2_n_166 & sub_613_2_n_88));
 assign sub_613_2_n_168 = ~(sub_613_2_n_80 | (sub_613_2_n_165 & sub_613_2_n_73));
 assign sub_613_2_n_167 = ~(sub_613_2_n_162 & sub_613_2_n_130);
 assign sub_613_2_n_166 = ~(sub_613_2_n_146 & (sub_613_2_n_160 | sub_613_2_n_136));
 assign sub_613_2_n_165 = ~(sub_613_2_n_125 & (sub_613_2_n_160 | sub_613_2_n_107));
 assign sub_613_2_n_164 = ~(sub_613_2_n_62 & (sub_613_2_n_160 | sub_613_2_n_2));
 assign in1_61_8_ = ~(sub_613_2_n_160 ^ sub_613_2_n_16);
 assign sub_613_2_n_162 = ~(sub_613_2_n_150 & (sub_613_2_n_160 | sub_613_2_n_140));
 assign sub_613_2_n_161 = ~(sub_613_2_n_70 | ~(sub_613_2_n_158 | sub_613_2_n_15));
 assign sub_613_2_n_160 = ~(sub_613_2_n_159 | sub_613_2_n_144);
 assign sub_613_2_n_159 = ~(sub_613_2_n_154 | (sub_613_2_n_17 | sub_613_2_n_20));
 assign sub_613_2_n_158 = ~(sub_613_2_n_138 | (sub_613_2_n_155 & sub_613_2_n_120));
 assign sub_613_2_n_157 = ~(sub_613_2_n_84 | (sub_613_2_n_155 & sub_613_2_n_14));
 assign in1_61_2_ = ~(sub_613_2_n_153 & ~sub_613_2_n_152);
 assign sub_613_2_n_155 = ~sub_613_2_n_154;
 assign sub_613_2_n_154 = ~(sub_613_2_n_151 | sub_613_2_n_124);
 assign sub_613_2_n_153 = ~(sub_613_2_n_148 & sub_613_2_n_98);
 assign sub_613_2_n_152 = ~(sub_613_2_n_148 | sub_613_2_n_98);
 assign sub_613_2_n_151 = ~(sub_613_2_n_142 | sub_613_2_n_111);
 assign sub_613_2_n_150 = ~(sub_613_2_n_147 | sub_613_2_n_145);
 assign sub_613_2_n_149 = ~(sub_613_2_n_131 & (sub_613_2_n_143 | sub_613_2_n_132));
 assign sub_613_2_n_148 = ~sub_613_2_n_142;
 assign sub_613_2_n_147 = ~(sub_613_2_n_146 | sub_613_2_n_134);
 assign sub_613_2_n_146 = ~(sub_613_2_n_37 | sub_613_2_n_129);
 assign sub_613_2_n_145 = ~(sub_613_2_n_121 & (sub_613_2_n_128 | sub_613_2_n_18));
 assign sub_613_2_n_144 = ~(sub_613_2_n_122 & (sub_613_2_n_137 | sub_613_2_n_20));
 assign sub_613_2_n_143 = ~(sub_613_2_n_31 | sub_613_2_n_123);
 assign sub_613_2_n_142 = ~(sub_613_2_n_141 | sub_613_2_n_78);
 assign sub_613_2_n_141 = ~(sub_613_2_n_139 | ~(in1_59_0_ | sub_613_2_n_59));
 assign sub_613_2_n_140 = ~(sub_613_2_n_135 & sub_613_2_n_133);
 assign sub_613_2_n_139 = ~sub_613_2_n_61;
 assign sub_613_2_n_138 = ~sub_613_2_n_137;
 assign sub_613_2_n_136 = ~sub_613_2_n_135;
 assign sub_613_2_n_134 = ~sub_613_2_n_133;
 assign sub_613_2_n_131 = ~(in1_59_19_ & (sub_613_2_n_97 & ~{in2[20]}));
 assign sub_613_2_n_130 = (sub_613_2_n_116 & sub_613_2_n_104);
 assign sub_613_2_n_129 = ~(sub_613_2_n_90 & (sub_613_2_n_79 | sub_613_2_n_0));
 assign sub_613_2_n_137 = ~(sub_613_2_n_96 | sub_613_2_n_8);
 assign sub_613_2_n_135 = (sub_613_2_n_106 & sub_613_2_n_118);
 assign sub_613_2_n_133 = ~(sub_613_2_n_18 | ~sub_613_2_n_113);
 assign sub_613_2_n_132 = ~(sub_613_2_n_97 & sub_613_2_n_1);
 assign sub_613_2_n_127 = ~sub_613_2_n_126;
 assign sub_613_2_n_124 = ~(sub_613_2_n_91 & (sub_613_2_n_87 | sub_613_2_n_5));
 assign sub_613_2_n_123 = ~(sub_613_2_n_92 & (sub_613_2_n_66 | sub_613_2_n_3));
 assign sub_613_2_n_122 = ~(sub_613_2_n_12 | ~(sub_613_2_n_69 | sub_613_2_n_48));
 assign sub_613_2_n_121 = ~(sub_613_2_n_9 | ~(sub_613_2_n_71 | sub_613_2_n_75));
 assign sub_613_2_n_128 = ~(sub_613_2_n_110 | sub_613_2_n_10);
 assign sub_613_2_n_126 = ~(sub_613_2_n_112 | sub_613_2_n_76);
 assign sub_613_2_n_125 = ~(sub_613_2_n_95 | sub_613_2_n_4);
 assign sub_613_2_n_120 = ~sub_613_2_n_17;
 assign sub_613_2_n_115 = ~sub_613_2_n_114;
 assign sub_613_2_n_112 = ~(sub_613_2_n_85 | sub_613_2_n_81);
 assign sub_613_2_n_111 = ~(sub_613_2_n_89 & ~sub_613_2_n_74);
 assign sub_613_2_n_110 = ~(sub_613_2_n_64 | sub_613_2_n_82);
 assign sub_613_2_n_119 = ~(sub_613_2_n_70 | sub_613_2_n_15);
 assign sub_613_2_n_118 = ~(sub_613_2_n_45 | sub_613_2_n_0);
 assign sub_613_2_n_117 = ~(sub_613_2_n_76 | sub_613_2_n_81);
 assign sub_613_2_n_116 = ~(sub_613_2_n_6 | sub_613_2_n_81);
 assign sub_613_2_n_109 = ~(sub_613_2_n_85 & sub_613_2_n_63);
 assign sub_613_2_n_114 = ~(sub_613_2_n_9 | sub_613_2_n_75);
 assign sub_613_2_n_113 = ~(sub_613_2_n_7 | sub_613_2_n_82);
 assign sub_613_2_n_107 = ~sub_613_2_n_106;
 assign sub_613_2_n_96 = ~(sub_613_2_n_83 | sub_613_2_n_47);
 assign sub_613_2_n_95 = ~(sub_613_2_n_62 | sub_613_2_n_68);
 assign in1_61_0_ = ~(sub_613_2_n_61 & ~(sub_613_2_n_50 & {in1[28]}));
 assign sub_613_2_n_108 = ~(sub_613_2_n_10 | sub_613_2_n_82);
 assign sub_613_2_n_106 = ~(sub_613_2_n_2 | sub_613_2_n_68);
 assign sub_613_2_n_105 = ~(sub_613_2_n_80 | sub_613_2_n_45);
 assign sub_613_2_n_104 = ~(sub_613_2_n_13 | sub_613_2_n_3);
 assign sub_613_2_n_103 = ~(sub_613_2_n_4 | sub_613_2_n_68);
 assign sub_613_2_n_102 = ~(sub_613_2_n_12 | sub_613_2_n_48);
 assign sub_613_2_n_101 = ~(sub_613_2_n_65 | sub_613_2_n_7);
 assign sub_613_2_n_100 = ~(sub_613_2_n_8 | sub_613_2_n_47);
 assign sub_613_2_n_99 = ~(sub_613_2_n_72 | sub_613_2_n_46);
 assign sub_613_2_n_98 = ~(sub_613_2_n_87 & ~sub_613_2_n_74);
 assign sub_613_2_n_97 = ~({in2[22]} | ({in2[23]} | {in2[21]}));
 assign sub_613_2_n_93 = ~(sub_613_2_n_67 | sub_613_2_n_13);
 assign sub_613_2_n_89 = ~sub_613_2_n_5;
 assign sub_613_2_n_88 = ~sub_613_2_n_7;
 assign sub_613_2_n_86 = ~sub_613_2_n_85;
 assign sub_613_2_n_84 = ~sub_613_2_n_83;
 assign sub_613_2_n_80 = ~sub_613_2_n_79;
 assign sub_613_2_n_92 = ~(in1_59_18_ & ~{in2[19]});
 assign sub_613_2_n_91 = ~(in1_59_2_ & ~{in2[3]});
 assign sub_613_2_n_90 = ~(in1_59_10_ & ~{in2[11]});
 assign sub_613_2_n_78 = ~(sub_613_2_n_58 | ~sub_613_2_n_59);
 assign sub_613_2_n_77 = ~({in2[20]} | ~in1_59_19_);
 assign sub_613_2_n_87 = ~(in1_59_1_ & ~{in2[2]});
 assign sub_613_2_n_85 = ~(in1_59_15_ & ~{in2[16]});
 assign sub_613_2_n_83 = ~(in1_59_3_ & ~{in2[4]});
 assign sub_613_2_n_82 = ~(in1_59_12_ | sub_613_2_n_57);
 assign sub_613_2_n_81 = ~(in1_59_16_ | sub_613_2_n_53);
 assign sub_613_2_n_79 = ~(in1_59_9_ & ~{in2[10]});
 assign sub_613_2_n_48 = ~(in1_59_6_ | sub_613_2_n_60);
 assign sub_613_2_n_73 = ~sub_613_2_n_45;
 assign sub_613_2_n_72 = ~sub_613_2_n_71;
 assign sub_613_2_n_70 = ~sub_613_2_n_69;
 assign sub_613_2_n_67 = ~sub_613_2_n_66;
 assign sub_613_2_n_65 = ~sub_613_2_n_64;
 assign sub_613_2_n_63 = ~sub_613_2_n_6;
 assign sub_613_2_n_76 = (sub_613_2_n_53 & in1_59_16_);
 assign sub_613_2_n_75 = ~(in1_59_14_ | sub_613_2_n_51);
 assign sub_613_2_n_74 = ~(in1_59_1_ | ~{in2[2]});
 assign sub_613_2_n_71 = ~(in1_59_13_ & ~{in2[14]});
 assign sub_613_2_n_69 = ~(in1_59_5_ & ~{in2[6]});
 assign sub_613_2_n_47 = ~(in1_59_4_ | sub_613_2_n_55);
 assign sub_613_2_n_68 = ~(in1_59_8_ | sub_613_2_n_54);
 assign sub_613_2_n_66 = ~(in1_59_17_ & ~{in2[18]});
 assign sub_613_2_n_64 = ~(in1_59_11_ & ~{in2[12]});
 assign sub_613_2_n_62 = ~(in1_59_7_ & ~{in2[8]});
 assign sub_613_2_n_61 = ~({in2[0]} & ~{in1[28]});
 assign sub_613_2_n_60 = ~{in2[7]};
 assign sub_613_2_n_59 = ~{in2[1]};
 assign sub_613_2_n_58 = ~in1_59_0_;
 assign sub_613_2_n_57 = ~{in2[13]};
 assign sub_613_2_n_56 = ~{in2[10]};
 assign sub_613_2_n_55 = ~{in2[5]};
 assign sub_613_2_n_54 = ~{in2[9]};
 assign sub_613_2_n_53 = ~{in2[17]};
 assign sub_613_2_n_52 = ~{in2[14]};
 assign sub_613_2_n_51 = ~{in2[15]};
 assign sub_613_2_n_50 = ~{in2[0]};
 assign sub_613_2_n_46 = ~(in1_59_13_ | sub_613_2_n_52);
 assign sub_613_2_n_45 = ~(in1_59_9_ | sub_613_2_n_56);
 assign sub_613_2_n_44 = ~(sub_613_2_n_72 | ~(sub_613_2_n_40 | sub_613_2_n_46));
 assign sub_613_2_n_43 = (sub_613_2_n_167 & sub_613_2_n_143);
 assign sub_613_2_n_42 = (sub_613_2_n_166 & sub_613_2_n_113);
 assign in1_61_4_ = (sub_613_2_n_155 ^ sub_613_2_n_21);
 assign sub_613_2_n_40 = ~(sub_613_2_n_42 | ~sub_613_2_n_128);
 assign in1_61_6_ = ~(sub_613_2_n_158 ^ sub_613_2_n_119);
 assign in1_61_3_ = ~(sub_613_2_n_22 ^ sub_613_2_n_25);
 assign sub_613_2_n_37 = ~(sub_613_2_n_125 | ~sub_613_2_n_118);
 assign in1_61_20_ = ~(sub_613_2_n_43 ^ sub_613_2_n_19);
 assign in1_61_17_ = ~(sub_613_2_n_171 ^ sub_613_2_n_117);
 assign in1_61_13_ = ~(sub_613_2_n_169 ^ sub_613_2_n_108);
 assign in1_61_11_ = ~(sub_613_2_n_168 ^ sub_613_2_n_24);
 assign in1_61_10_ = (sub_613_2_n_165 ^ sub_613_2_n_105);
 assign sub_613_2_n_31 = ~(sub_613_2_n_126 | ~sub_613_2_n_104);
 assign in1_61_9_ = (sub_613_2_n_164 ^ sub_613_2_n_103);
 assign in1_61_7_ = ~(sub_613_2_n_161 ^ sub_613_2_n_102);
 assign in1_61_12_ = (sub_613_2_n_166 ^ sub_613_2_n_101);
 assign in1_61_5_ = ~(sub_613_2_n_157 ^ sub_613_2_n_100);
 assign in1_61_14_ = ~(sub_613_2_n_40 ^ sub_613_2_n_99);
 assign sub_613_2_n_25 = ~(sub_613_2_n_5 | ~sub_613_2_n_91);
 assign sub_613_2_n_24 = ~(sub_613_2_n_0 | ~sub_613_2_n_90);
 assign sub_613_2_n_23 = ~(sub_613_2_n_92 & ~sub_613_2_n_3);
 assign sub_613_2_n_22 = (sub_613_2_n_87 & (sub_613_2_n_142 | sub_613_2_n_74));
 assign sub_613_2_n_21 = ~(sub_613_2_n_84 | ~sub_613_2_n_14);
 assign sub_613_2_n_20 = (sub_613_2_n_48 | sub_613_2_n_15);
 assign sub_613_2_n_19 = ~(sub_613_2_n_77 | ~sub_613_2_n_1);
 assign sub_613_2_n_18 = (sub_613_2_n_75 | sub_613_2_n_46);
 assign sub_613_2_n_17 = ~(sub_613_2_n_14 & ~sub_613_2_n_47);
 assign sub_613_2_n_16 = ~(sub_613_2_n_2 | ~sub_613_2_n_62);
 assign sub_613_2_n_15 = ~(in1_59_5_ | ~{in2[6]});
 assign sub_613_2_n_14 = ~({in2[4]} & ~in1_59_3_);
 assign sub_613_2_n_13 = ~(in1_59_17_ | ~{in2[18]});
 assign sub_613_2_n_12 = (in1_59_6_ & sub_613_2_n_60);
 assign sub_613_2_n_10 = (in1_59_12_ & sub_613_2_n_57);
 assign sub_613_2_n_9 = (in1_59_14_ & sub_613_2_n_51);
 assign sub_613_2_n_8 = (in1_59_4_ & sub_613_2_n_55);
 assign sub_613_2_n_7 = ~(in1_59_11_ | ~{in2[12]});
 assign sub_613_2_n_6 = ~(in1_59_15_ | ~{in2[16]});
 assign sub_613_2_n_5 = ~(in1_59_2_ | ~{in2[3]});
 assign sub_613_2_n_4 = (in1_59_8_ & sub_613_2_n_54);
 assign sub_613_2_n_3 = ~(in1_59_18_ | ~{in2[19]});
 assign sub_613_2_n_2 = ~(in1_59_7_ | ~{in2[8]});
 assign sub_613_2_n_1 = ~({in2[20]} & ~in1_59_19_);
 assign sub_613_2_n_0 = ~(in1_59_10_ | ~{in2[11]});
 assign in1_61_1_ = (sub_613_2_n_58 ^ ({in2[1]} ^ sub_613_2_n_61));
 assign in1_64_21_ = (n_1518 ^ n_1520);
 assign in1_64_19_ = ~((sub_634_2_n_113 & ~sub_634_2_n_167) | (sub_634_2_n_112 & sub_634_2_n_167));
 assign sub_634_2_n_168 = ~(sub_634_2_n_70 | (sub_634_2_n_161 & sub_634_2_n_9));
 assign sub_634_2_n_167 = ~(sub_634_2_n_67 & (sub_634_2_n_160 | sub_634_2_n_14));
 assign in1_64_17_ = ~(sub_634_2_n_159 ^ sub_634_2_n_18);
 assign sub_634_2_n_165 = ~(sub_634_2_n_64 & (sub_634_2_n_156 | sub_634_2_n_65));
 assign in1_64_14_ = ~(sub_634_2_n_155 ^ sub_634_2_n_91);
 assign in1_64_13_ = ~(sub_634_2_n_154 ^ sub_634_2_n_93);
 assign in1_64_11_ = ~(sub_634_2_n_153 ^ sub_634_2_n_92);
 assign sub_634_2_n_161 = ~(sub_634_2_n_132 & (sub_634_2_n_49 | sub_634_2_n_124));
 assign sub_634_2_n_160 = ~(sub_634_2_n_38 | sub_634_2_n_125);
 assign sub_634_2_n_159 = ~(sub_634_2_n_81 & (sub_634_2_n_49 | sub_634_2_n_66));
 assign in1_64_24_ = ~(sub_634_2_n_157 | sub_634_2_n_137);
 assign sub_634_2_n_157 = ~(sub_634_2_n_151 | sub_634_2_n_44);
 assign sub_634_2_n_156 = ~sub_634_2_n_155;
 assign sub_634_2_n_155 = ~(sub_634_2_n_118 & (sub_634_2_n_46 | sub_634_2_n_108));
 assign sub_634_2_n_154 = ~(sub_634_2_n_82 & (sub_634_2_n_46 | sub_634_2_n_12));
 assign sub_634_2_n_153 = ~(sub_634_2_n_83 & (sub_634_2_n_149 | sub_634_2_n_85));
 assign in1_64_12_ = ~(sub_634_2_n_46 ^ sub_634_2_n_27);
 assign sub_634_2_n_151 = ~(sub_634_2_n_150 | sub_634_2_n_138);
 assign sub_634_2_n_150 = ~(sub_634_2_n_144 | (sub_634_2_n_40 | sub_634_2_n_32));
 assign sub_634_2_n_149 = ~sub_634_2_n_148;
 assign sub_634_2_n_148 = ~(sub_634_2_n_119 & (sub_634_2_n_144 | sub_634_2_n_99));
 assign sub_634_2_n_147 = ~(sub_634_2_n_63 & (sub_634_2_n_144 | sub_634_2_n_10));
 assign sub_634_2_n_146 = ~(sub_634_2_n_144 | sub_634_2_n_40);
 assign sub_634_2_n_145 = ~(sub_634_2_n_71 & (sub_634_2_n_43 | sub_634_2_n_5));
 assign sub_634_2_n_144 = ~(sub_634_2_n_143 | sub_634_2_n_130);
 assign sub_634_2_n_143 = ~(sub_634_2_n_140 | (sub_634_2_n_16 | sub_634_2_n_20));
 assign sub_634_2_n_142 = ~(sub_634_2_n_80 & (sub_634_2_n_140 | sub_634_2_n_68));
 assign sub_634_2_n_141 = ~(sub_634_2_n_52 & (sub_634_2_n_136 | sub_634_2_n_7));
 assign sub_634_2_n_140 = ~(sub_634_2_n_139 | sub_634_2_n_121);
 assign sub_634_2_n_139 = ~(sub_634_2_n_136 | sub_634_2_n_28);
 assign sub_634_2_n_138 = ~(sub_634_2_n_131 & (sub_634_2_n_133 | sub_634_2_n_32));
 assign sub_634_2_n_137 = ~(sub_634_2_n_128 & (sub_634_2_n_132 | sub_634_2_n_122));
 assign sub_634_2_n_136 = ~(sub_634_2_n_135 | sub_634_2_n_62);
 assign sub_634_2_n_135 = ~(sub_634_2_n_129 & sub_634_2_n_45);
 assign in1_64_1_ = ~(in1_62_0_ ^ ({in2[1]} ^ sub_634_2_n_77));
 assign sub_634_2_n_133 = ~(sub_634_2_n_127 | sub_634_2_n_114);
 assign sub_634_2_n_132 = ~(sub_634_2_n_115 | (sub_634_2_n_125 & sub_634_2_n_102));
 assign sub_634_2_n_131 = ~(sub_634_2_n_126 | sub_634_2_n_116);
 assign sub_634_2_n_130 = ~(sub_634_2_n_117 & (sub_634_2_n_120 | sub_634_2_n_20));
 assign sub_634_2_n_129 = ~(sub_634_2_n_77 & ~{in2[1]});
 assign sub_634_2_n_128 = ~(sub_634_2_n_89 & (sub_634_2_n_94 | sub_634_2_n_75));
 assign sub_634_2_n_127 = ~(sub_634_2_n_110 | sub_634_2_n_119);
 assign sub_634_2_n_126 = ~(sub_634_2_n_118 | sub_634_2_n_15);
 assign sub_634_2_n_124 = ~sub_634_2_n_123;
 assign sub_634_2_n_121 = ~(sub_634_2_n_74 & (sub_634_2_n_52 | sub_634_2_n_4));
 assign sub_634_2_n_125 = ~(sub_634_2_n_90 & (sub_634_2_n_81 | sub_634_2_n_3));
 assign sub_634_2_n_123 = (sub_634_2_n_109 & sub_634_2_n_102);
 assign sub_634_2_n_122 = ~(sub_634_2_n_105 & sub_634_2_n_9);
 assign sub_634_2_n_117 = ~(sub_634_2_n_97 | sub_634_2_n_87);
 assign sub_634_2_n_116 = ~(sub_634_2_n_73 & (sub_634_2_n_64 | sub_634_2_n_6));
 assign sub_634_2_n_115 = ~(sub_634_2_n_76 & (sub_634_2_n_67 | sub_634_2_n_13));
 assign sub_634_2_n_114 = ~(sub_634_2_n_104 & sub_634_2_n_86);
 assign sub_634_2_n_120 = ~(sub_634_2_n_95 | sub_634_2_n_8);
 assign sub_634_2_n_119 = ~(sub_634_2_n_106 | sub_634_2_n_0);
 assign sub_634_2_n_118 = ~(sub_634_2_n_88 | ~(sub_634_2_n_82 | sub_634_2_n_84));
 assign sub_634_2_n_113 = ~sub_634_2_n_112;
 assign sub_634_2_n_108 = ~sub_634_2_n_107;
 assign sub_634_2_n_106 = ~(sub_634_2_n_63 | sub_634_2_n_79);
 assign sub_634_2_n_105 = ~(sub_634_2_n_78 | ~sub_634_2_n_89);
 assign sub_634_2_n_104 = ~(sub_634_2_n_72 & ~sub_634_2_n_83);
 assign sub_634_2_n_103 = ~(sub_634_2_n_69 & sub_634_2_n_9);
 assign sub_634_2_n_112 = ~(sub_634_2_n_13 | ~sub_634_2_n_76);
 assign sub_634_2_n_111 = ~(sub_634_2_n_87 | sub_634_2_n_51);
 assign sub_634_2_n_110 = ~(sub_634_2_n_72 & ~sub_634_2_n_85);
 assign sub_634_2_n_109 = ~(sub_634_2_n_66 | sub_634_2_n_3);
 assign sub_634_2_n_107 = ~(sub_634_2_n_12 | sub_634_2_n_84);
 assign sub_634_2_n_99 = ~sub_634_2_n_98;
 assign sub_634_2_n_97 = ~(sub_634_2_n_71 | sub_634_2_n_51);
 assign in1_64_0_ = ~(sub_634_2_n_77 & ~(sub_634_2_n_59 & {in1[27]}));
 assign sub_634_2_n_95 = ~(sub_634_2_n_80 | sub_634_2_n_50);
 assign sub_634_2_n_94 = ~(sub_634_2_n_69 | sub_634_2_n_78);
 assign sub_634_2_n_93 = (sub_634_2_n_88 | sub_634_2_n_84);
 assign sub_634_2_n_92 = ~(sub_634_2_n_86 & sub_634_2_n_72);
 assign sub_634_2_n_102 = ~(sub_634_2_n_14 | sub_634_2_n_13);
 assign sub_634_2_n_91 = ~(sub_634_2_n_64 & ~sub_634_2_n_65);
 assign sub_634_2_n_101 = ~(sub_634_2_n_0 | sub_634_2_n_79);
 assign sub_634_2_n_100 = ~(sub_634_2_n_8 | sub_634_2_n_50);
 assign sub_634_2_n_98 = ~(sub_634_2_n_10 | sub_634_2_n_79);
 assign sub_634_2_n_90 = ~(in1_62_16_ & ~{in2[17]});
 assign sub_634_2_n_89 = ~({in2[22]} | {in2[23]});
 assign sub_634_2_n_88 = (sub_634_2_n_57 & in1_62_12_);
 assign sub_634_2_n_87 = (sub_634_2_n_55 & in1_62_6_);
 assign sub_634_2_n_86 = ~(in1_62_10_ & ~{in2[11]});
 assign sub_634_2_n_85 = ~(in1_62_9_ | ~{in2[10]});
 assign sub_634_2_n_84 = ~(in1_62_12_ | sub_634_2_n_57);
 assign sub_634_2_n_83 = ~(in1_62_9_ & ~{in2[10]});
 assign sub_634_2_n_82 = ~(in1_62_11_ & ~{in2[12]});
 assign sub_634_2_n_81 = ~(in1_62_15_ & ~{in2[16]});
 assign sub_634_2_n_52 = ~(in1_62_1_ & ~{in2[2]});
 assign sub_634_2_n_80 = ~(in1_62_3_ & ~{in2[4]});
 assign sub_634_2_n_79 = ~(in1_62_8_ | sub_634_2_n_56);
 assign sub_634_2_n_78 = ~(in1_62_20_ | sub_634_2_n_60);
 assign sub_634_2_n_77 = ~({in2[0]} & ~{in1[27]});
 assign sub_634_2_n_70 = ~sub_634_2_n_69;
 assign sub_634_2_n_68 = ~sub_634_2_n_11;
 assign sub_634_2_n_76 = ~(in1_62_18_ & ~{in2[19]});
 assign sub_634_2_n_75 = (sub_634_2_n_60 & in1_62_20_);
 assign sub_634_2_n_74 = ~(in1_62_2_ & ~{in2[3]});
 assign sub_634_2_n_73 = ~(in1_62_14_ & ~{in2[15]});
 assign sub_634_2_n_62 = (sub_634_2_n_54 & in1_62_0_);
 assign sub_634_2_n_72 = ~(sub_634_2_n_58 & {in2[11]});
 assign sub_634_2_n_51 = ~(in1_62_6_ | sub_634_2_n_55);
 assign sub_634_2_n_71 = ~(in1_62_5_ & ~{in2[6]});
 assign sub_634_2_n_69 = ~(in1_62_19_ & ~{in2[20]});
 assign sub_634_2_n_67 = ~(in1_62_17_ & ~{in2[18]});
 assign sub_634_2_n_66 = ~(in1_62_15_ | ~{in2[16]});
 assign sub_634_2_n_65 = ~(in1_62_13_ | ~{in2[14]});
 assign sub_634_2_n_50 = ~(in1_62_4_ | sub_634_2_n_61);
 assign sub_634_2_n_64 = ~(in1_62_13_ & ~{in2[14]});
 assign sub_634_2_n_63 = ~(in1_62_7_ & ~{in2[8]});
 assign sub_634_2_n_61 = ~{in2[5]};
 assign sub_634_2_n_60 = ~{in2[21]};
 assign sub_634_2_n_59 = ~{in2[0]};
 assign sub_634_2_n_58 = ~in1_62_10_;
 assign sub_634_2_n_57 = ~{in2[13]};
 assign sub_634_2_n_56 = ~{in2[9]};
 assign sub_634_2_n_55 = ~{in2[7]};
 assign sub_634_2_n_54 = ~{in2[1]};
 assign sub_634_2_n_49 = sub_634_2_n_151;
 assign in1_64_20_ = ~(sub_634_2_n_161 ^ sub_634_2_n_103);
 assign in1_64_18_ = ~(sub_634_2_n_160 ^ sub_634_2_n_17);
 assign sub_634_2_n_46 = ~(sub_634_2_n_146 | ~sub_634_2_n_133);
 assign sub_634_2_n_45 = ~(in1_62_0_ & sub_634_2_n_77);
 assign sub_634_2_n_44 = ~(sub_634_2_n_123 & ~sub_634_2_n_122);
 assign sub_634_2_n_43 = (sub_634_2_n_120 & (sub_634_2_n_140 | sub_634_2_n_16));
 assign in1_64_7_ = (sub_634_2_n_145 ^ sub_634_2_n_111);
 assign in1_64_3_ = (sub_634_2_n_141 ^ sub_634_2_n_22);
 assign sub_634_2_n_40 = ~(sub_634_2_n_98 & ~sub_634_2_n_110);
 assign in1_64_2_ = ~(sub_634_2_n_136 ^ sub_634_2_n_25);
 assign sub_634_2_n_38 = ~(sub_634_2_n_49 | ~sub_634_2_n_109);
 assign in1_64_8_ = ~(sub_634_2_n_144 ^ sub_634_2_n_2);
 assign in1_64_4_ = ~(sub_634_2_n_140 ^ sub_634_2_n_24);
 assign in1_64_6_ = ~(sub_634_2_n_43 ^ sub_634_2_n_19);
 assign in1_64_10_ = (sub_634_2_n_148 ^ sub_634_2_n_1);
 assign in1_64_9_ = (sub_634_2_n_147 ^ sub_634_2_n_101);
 assign sub_634_2_n_32 = ~(sub_634_2_n_107 & ~sub_634_2_n_15);
 assign in1_64_5_ = (sub_634_2_n_142 ^ sub_634_2_n_100);
 assign in1_64_16_ = ~(sub_634_2_n_49 ^ sub_634_2_n_26);
 assign in1_64_15_ = (sub_634_2_n_165 ^ sub_634_2_n_21);
 assign sub_634_2_n_28 = (sub_634_2_n_4 | sub_634_2_n_7);
 assign sub_634_2_n_27 = ~(sub_634_2_n_12 | ~sub_634_2_n_82);
 assign sub_634_2_n_26 = ~(sub_634_2_n_66 | ~sub_634_2_n_81);
 assign sub_634_2_n_25 = ~(sub_634_2_n_7 | ~sub_634_2_n_52);
 assign sub_634_2_n_24 = ~(sub_634_2_n_68 | ~sub_634_2_n_80);
 assign sub_634_2_n_23 = (sub_634_2_n_75 | sub_634_2_n_78);
 assign sub_634_2_n_22 = ~(sub_634_2_n_4 | ~sub_634_2_n_74);
 assign sub_634_2_n_21 = ~(sub_634_2_n_6 | ~sub_634_2_n_73);
 assign sub_634_2_n_20 = (sub_634_2_n_51 | sub_634_2_n_5);
 assign sub_634_2_n_19 = ~(sub_634_2_n_5 | ~sub_634_2_n_71);
 assign sub_634_2_n_18 = ~(sub_634_2_n_90 & ~sub_634_2_n_3);
 assign sub_634_2_n_17 = ~(sub_634_2_n_14 | ~sub_634_2_n_67);
 assign sub_634_2_n_16 = ~(sub_634_2_n_11 & ~sub_634_2_n_50);
 assign sub_634_2_n_15 = (sub_634_2_n_6 | sub_634_2_n_65);
 assign sub_634_2_n_14 = ~(in1_62_17_ | ~{in2[18]});
 assign sub_634_2_n_13 = ~(in1_62_18_ | ~{in2[19]});
 assign sub_634_2_n_12 = ~(in1_62_11_ | ~{in2[12]});
 assign sub_634_2_n_11 = ~({in2[4]} & ~in1_62_3_);
 assign sub_634_2_n_10 = ~(in1_62_7_ | ~{in2[8]});
 assign sub_634_2_n_9 = ~({in2[20]} & ~in1_62_19_);
 assign sub_634_2_n_8 = (in1_62_4_ & sub_634_2_n_61);
 assign sub_634_2_n_7 = ~(in1_62_1_ | ~{in2[2]});
 assign sub_634_2_n_6 = ~(in1_62_14_ | ~{in2[15]});
 assign sub_634_2_n_5 = ~(in1_62_5_ | ~{in2[6]});
 assign sub_634_2_n_4 = ~(in1_62_2_ | ~{in2[3]});
 assign sub_634_2_n_3 = ~(in1_62_16_ | ~{in2[17]});
 assign sub_634_2_n_2 = ~(sub_634_2_n_10 | ~sub_634_2_n_63);
 assign sub_634_2_n_1 = ~(sub_634_2_n_85 | ~sub_634_2_n_83);
 assign sub_634_2_n_0 = (in1_62_8_ & sub_634_2_n_56);
 assign in1_67_22_ = ~(sub_655_2_n_178 ^ sub_655_2_n_114);
 assign in1_67_19_ = ~(sub_655_2_n_176 ^ sub_655_2_n_112);
 assign sub_655_2_n_178 = ~(sub_655_2_n_128 & (sub_655_2_n_49 | sub_655_2_n_106));
 assign sub_655_2_n_177 = ~(sub_655_2_n_69 & (sub_655_2_n_49 | sub_655_2_n_8));
 assign sub_655_2_n_176 = ~(sub_655_2_n_71 & (sub_655_2_n_43 | sub_655_2_n_4));
 assign in1_67_20_ = ~(sub_655_2_n_49 ^ sub_655_2_n_18);
 assign in1_67_24_ = ~(sub_655_2_n_171 | sub_655_2_n_147);
 assign sub_655_2_n_173 = ~(sub_655_2_n_75 & (sub_655_2_n_166 | sub_655_2_n_1));
 assign in1_67_14_ = ~(sub_655_2_n_165 ^ sub_655_2_n_97);
 assign sub_655_2_n_171 = ~(sub_655_2_n_167 | sub_655_2_n_132);
 assign sub_655_2_n_170 = ~(sub_655_2_n_89 & (sub_655_2_n_161 | sub_655_2_n_14));
 assign in1_67_16_ = ~(sub_655_2_n_161 ^ sub_655_2_n_25);
 assign sub_655_2_n_168 = ~(sub_655_2_n_161 | ~sub_655_2_n_109);
 assign sub_655_2_n_167 = ~(sub_655_2_n_160 & sub_655_2_n_41);
 assign sub_655_2_n_166 = ~sub_655_2_n_165;
 assign sub_655_2_n_165 = ~(sub_655_2_n_129 & (sub_655_2_n_45 | sub_655_2_n_121));
 assign sub_655_2_n_164 = ~(sub_655_2_n_77 & (sub_655_2_n_45 | sub_655_2_n_7));
 assign sub_655_2_n_163 = ~(sub_655_2_n_84 | (sub_655_2_n_159 & sub_655_2_n_88));
 assign in1_67_7_ = (sub_655_2_n_156 ^ sub_655_2_n_95);
 assign sub_655_2_n_161 = ~sub_655_2_n_160;
 assign sub_655_2_n_160 = ~(sub_655_2_n_148 & (sub_655_2_n_155 | (sub_655_2_n_37 | sub_655_2_n_135)));
 assign sub_655_2_n_159 = ~(sub_655_2_n_133 & (sub_655_2_n_155 | sub_655_2_n_108));
 assign sub_655_2_n_158 = ~(sub_655_2_n_68 & (sub_655_2_n_155 | sub_655_2_n_15));
 assign in1_67_8_ = ~(sub_655_2_n_155 ^ sub_655_2_n_17);
 assign sub_655_2_n_156 = ~(sub_655_2_n_72 & (sub_655_2_n_47 | sub_655_2_n_2));
 assign sub_655_2_n_155 = ~(sub_655_2_n_154 | sub_655_2_n_138);
 assign sub_655_2_n_154 = ~(sub_655_2_n_53 | (sub_655_2_n_27 | sub_655_2_n_22));
 assign sub_655_2_n_153 = ~(sub_655_2_n_67 & (sub_655_2_n_53 | sub_655_2_n_85));
 assign in1_67_2_ = ~(sub_655_2_n_150 & ~sub_655_2_n_151);
 assign sub_655_2_n_53 = ~(sub_655_2_n_149 | sub_655_2_n_124);
 assign sub_655_2_n_151 = ~(sub_655_2_n_144 | sub_655_2_n_119);
 assign sub_655_2_n_150 = ~(sub_655_2_n_144 & sub_655_2_n_119);
 assign sub_655_2_n_149 = ~(sub_655_2_n_144 | sub_655_2_n_26);
 assign sub_655_2_n_148 = ~(sub_655_2_n_145 | sub_655_2_n_139);
 assign sub_655_2_n_147 = ~(sub_655_2_n_146 & sub_655_2_n_142);
 assign sub_655_2_n_146 = ~(sub_655_2_n_140 & ~sub_655_2_n_132);
 assign sub_655_2_n_145 = ~(sub_655_2_n_141 | sub_655_2_n_135);
 assign sub_655_2_n_144 = ~(sub_655_2_n_143 | sub_655_2_n_64);
 assign sub_655_2_n_143 = ~(sub_655_2_n_137 & sub_655_2_n_44);
 assign sub_655_2_n_142 = ~(sub_655_2_n_116 | (sub_655_2_n_127 & sub_655_2_n_118));
 assign sub_655_2_n_141 = ~(sub_655_2_n_136 | sub_655_2_n_131);
 assign sub_655_2_n_140 = ~(sub_655_2_n_125 & (sub_655_2_n_134 | sub_655_2_n_20));
 assign sub_655_2_n_139 = ~(sub_655_2_n_123 & (sub_655_2_n_129 | sub_655_2_n_21));
 assign sub_655_2_n_138 = ~(sub_655_2_n_126 & (sub_655_2_n_130 | sub_655_2_n_22));
 assign sub_655_2_n_137 = ~(n_1545 & ~n_1586);
 assign sub_655_2_n_136 = ~(sub_655_2_n_133 | sub_655_2_n_24);
 assign sub_655_2_n_131 = ~(sub_655_2_n_90 & (sub_655_2_n_83 | sub_655_2_n_10));
 assign sub_655_2_n_135 = ~(sub_655_2_n_120 & sub_655_2_n_113);
 assign sub_655_2_n_134 = ~(sub_655_2_n_115 | sub_655_2_n_91);
 assign sub_655_2_n_133 = ~(sub_655_2_n_100 | sub_655_2_n_6);
 assign sub_655_2_n_132 = ~(sub_655_2_n_105 & sub_655_2_n_118);
 assign sub_655_2_n_128 = ~sub_655_2_n_127;
 assign sub_655_2_n_126 = ~(sub_655_2_n_80 | ~(sub_655_2_n_72 | sub_655_2_n_51));
 assign sub_655_2_n_125 = ~(sub_655_2_n_78 | ~(sub_655_2_n_71 | sub_655_2_n_73));
 assign sub_655_2_n_124 = ~(sub_655_2_n_94 & (sub_655_2_n_65 | sub_655_2_n_12));
 assign sub_655_2_n_123 = ~(sub_655_2_n_93 | ~(sub_655_2_n_75 | sub_655_2_n_74));
 assign sub_655_2_n_130 = ~(sub_655_2_n_99 | sub_655_2_n_9);
 assign sub_655_2_n_129 = ~(sub_655_2_n_117 | sub_655_2_n_92);
 assign sub_655_2_n_127 = ~(sub_655_2_n_79 & (sub_655_2_n_69 | sub_655_2_n_13));
 assign sub_655_2_n_121 = ~sub_655_2_n_120;
 assign sub_655_2_n_117 = ~(sub_655_2_n_77 | sub_655_2_n_87);
 assign sub_655_2_n_116 = ~(sub_655_2_n_81 | n_1403);
 assign sub_655_2_n_115 = ~(sub_655_2_n_89 | sub_655_2_n_86);
 assign sub_655_2_n_122 = ~(sub_655_2_n_9 | sub_655_2_n_52);
 assign sub_655_2_n_120 = ~(sub_655_2_n_7 | sub_655_2_n_87);
 assign sub_655_2_n_119 = ~(sub_655_2_n_66 | sub_655_2_n_70);
 assign sub_655_2_n_114 = ~(sub_655_2_n_81 & ~sub_655_2_n_5);
 assign sub_655_2_n_118 = ~(sub_655_2_n_5 | n_1403);
 assign sub_655_2_n_113 = ~(sub_655_2_n_1 | sub_655_2_n_74);
 assign sub_655_2_n_112 = (sub_655_2_n_78 | sub_655_2_n_73);
 assign sub_655_2_n_111 = ~(sub_655_2_n_71 & ~sub_655_2_n_4);
 assign sub_655_2_n_108 = ~sub_655_2_n_107;
 assign sub_655_2_n_106 = ~sub_655_2_n_105;
 assign sub_655_2_n_100 = ~(sub_655_2_n_68 | sub_655_2_n_76);
 assign sub_655_2_n_99 = ~(sub_655_2_n_67 | sub_655_2_n_52);
 assign in1_67_0_ = ~(n_1545 & ~(sub_655_2_n_56 & n_1583));
 assign sub_655_2_n_110 = ~(sub_655_2_n_93 | sub_655_2_n_74);
 assign sub_655_2_n_109 = ~(sub_655_2_n_14 | sub_655_2_n_86);
 assign sub_655_2_n_97 = ~(sub_655_2_n_75 & ~sub_655_2_n_1);
 assign sub_655_2_n_107 = ~(sub_655_2_n_15 | sub_655_2_n_76);
 assign sub_655_2_n_105 = ~(sub_655_2_n_8 | sub_655_2_n_13);
 assign sub_655_2_n_104 = ~(sub_655_2_n_84 | sub_655_2_n_3);
 assign sub_655_2_n_103 = ~(sub_655_2_n_6 | sub_655_2_n_76);
 assign sub_655_2_n_96 = ~(sub_655_2_n_77 & ~sub_655_2_n_7);
 assign sub_655_2_n_95 = ~(sub_655_2_n_80 | sub_655_2_n_51);
 assign sub_655_2_n_102 = ~(sub_655_2_n_92 | sub_655_2_n_87);
 assign sub_655_2_n_101 = ~(sub_655_2_n_91 | sub_655_2_n_86);
 assign sub_655_2_n_88 = ~sub_655_2_n_3;
 assign sub_655_2_n_85 = ~sub_655_2_n_11;
 assign sub_655_2_n_84 = ~sub_655_2_n_83;
 assign sub_655_2_n_94 = ~(n_1476 & ~n_1579);
 assign sub_655_2_n_93 = (sub_655_2_n_55 & n_1490);
 assign sub_655_2_n_92 = (sub_655_2_n_61 & n_1526);
 assign sub_655_2_n_91 = (sub_655_2_n_63 & n_1499);
 assign sub_655_2_n_90 = ~(n_1513 & ~n_1555);
 assign sub_655_2_n_52 = ~(n_1514 | sub_655_2_n_60);
 assign sub_655_2_n_89 = ~(in1_65_15_ & ~n_1549);
 assign sub_655_2_n_87 = ~(n_1526 | sub_655_2_n_61);
 assign sub_655_2_n_86 = ~(n_1499 | sub_655_2_n_63);
 assign sub_655_2_n_83 = ~(n_1504 & ~n_1551);
 assign sub_655_2_n_82 = ~({in2[0]} & ~{in1[26]});
 assign sub_655_2_n_66 = ~sub_655_2_n_65;
 assign sub_655_2_n_81 = ~(in1_65_21_ & ~n_1591);
 assign sub_655_2_n_80 = (sub_655_2_n_59 & n_1507);
 assign sub_655_2_n_79 = ~(in1_65_20_ & ~n_1593);
 assign sub_655_2_n_78 = (sub_655_2_n_57 & in1_65_18_);
 assign sub_655_2_n_64 = ~(sub_655_2_n_54 | ~sub_655_2_n_58);
 assign sub_655_2_n_77 = ~(n_1481 & ~n_1595);
 assign sub_655_2_n_51 = ~(n_1507 | sub_655_2_n_59);
 assign sub_655_2_n_76 = ~(n_1505 | sub_655_2_n_62);
 assign sub_655_2_n_75 = ~(n_1516 & ~n_1577);
 assign sub_655_2_n_74 = ~(n_1490 | sub_655_2_n_55);
 assign sub_655_2_n_73 = ~(in1_65_18_ | sub_655_2_n_57);
 assign sub_655_2_n_72 = ~(n_1508 & ~n_1567);
 assign sub_655_2_n_71 = ~(in1_65_17_ & ~n_1472);
 assign sub_655_2_n_70 = ~(n_1533 | ~n_1477);
 assign sub_655_2_n_69 = ~(in1_65_19_ & ~n_1565);
 assign sub_655_2_n_68 = ~(n_1506 & ~n_1479);
 assign sub_655_2_n_67 = ~(n_1515 & ~n_1535);
 assign sub_655_2_n_65 = ~(n_1533 & ~n_1477);
 assign sub_655_2_n_63 = ~n_1562;
 assign sub_655_2_n_62 = ~n_1589;
 assign sub_655_2_n_61 = ~n_1581;
 assign sub_655_2_n_60 = ~n_1569;
 assign sub_655_2_n_59 = ~n_1527;
 assign sub_655_2_n_58 = ~n_1586;
 assign sub_655_2_n_57 = ~n_1558;
 assign sub_655_2_n_56 = ~n_1543;
 assign sub_655_2_n_55 = ~n_1495;
 assign sub_655_2_n_54 = ~n_1529;
 assign in1_67_18_ = (sub_655_2_n_43 ^ sub_655_2_n_111);
 assign sub_655_2_n_49 = ~(sub_655_2_n_140 | ~sub_655_2_n_167);
 assign in1_67_12_ = (sub_655_2_n_45 ^ sub_655_2_n_96);
 assign sub_655_2_n_47 = (sub_655_2_n_130 & (sub_655_2_n_53 | sub_655_2_n_27));
 assign sub_655_2_n_46 = ~(sub_655_2_n_66 | ~(sub_655_2_n_144 | sub_655_2_n_70));
 assign sub_655_2_n_45 = (sub_655_2_n_141 & (sub_655_2_n_155 | sub_655_2_n_37));
 assign sub_655_2_n_44 = ~(n_1529 & n_1545);
 assign sub_655_2_n_43 = ~(sub_655_2_n_168 | ~sub_655_2_n_134);
 assign in1_67_5_ = (sub_655_2_n_153 ^ sub_655_2_n_122);
 assign sub_655_2_n_41 = ~(sub_655_2_n_20 | ~sub_655_2_n_109);
 assign in1_67_4_ = ~(sub_655_2_n_53 ^ sub_655_2_n_16);
 assign in1_67_21_ = (sub_655_2_n_177 ^ sub_655_2_n_23);
 assign in1_67_3_ = ~(sub_655_2_n_46 ^ sub_655_2_n_29);
 assign sub_655_2_n_37 = ~(sub_655_2_n_107 & ~sub_655_2_n_24);
 assign in1_67_15_ = (sub_655_2_n_173 ^ sub_655_2_n_110);
 assign in1_67_11_ = ~(sub_655_2_n_163 ^ sub_655_2_n_28);
 assign in1_67_10_ = (sub_655_2_n_159 ^ sub_655_2_n_104);
 assign in1_67_9_ = (sub_655_2_n_158 ^ sub_655_2_n_103);
 assign in1_67_6_ = ~(sub_655_2_n_47 ^ sub_655_2_n_19);
 assign in1_67_13_ = (sub_655_2_n_164 ^ sub_655_2_n_102);
 assign in1_67_17_ = (sub_655_2_n_170 ^ sub_655_2_n_101);
 assign sub_655_2_n_29 = ~(sub_655_2_n_12 | ~sub_655_2_n_94);
 assign sub_655_2_n_28 = ~(sub_655_2_n_10 | ~sub_655_2_n_90);
 assign sub_655_2_n_27 = ~(sub_655_2_n_11 & ~sub_655_2_n_52);
 assign sub_655_2_n_26 = (sub_655_2_n_12 | sub_655_2_n_70);
 assign sub_655_2_n_25 = ~(sub_655_2_n_14 | ~sub_655_2_n_89);
 assign sub_655_2_n_24 = (sub_655_2_n_10 | sub_655_2_n_3);
 assign sub_655_2_n_23 = ~(sub_655_2_n_13 | ~sub_655_2_n_79);
 assign sub_655_2_n_22 = (sub_655_2_n_51 | sub_655_2_n_2);
 assign sub_655_2_n_21 = (sub_655_2_n_74 | sub_655_2_n_1);
 assign sub_655_2_n_20 = (sub_655_2_n_73 | sub_655_2_n_4);
 assign sub_655_2_n_19 = ~(sub_655_2_n_2 | ~sub_655_2_n_72);
 assign sub_655_2_n_18 = ~(sub_655_2_n_8 | ~sub_655_2_n_69);
 assign sub_655_2_n_17 = ~(sub_655_2_n_15 | ~sub_655_2_n_68);
 assign sub_655_2_n_16 = ~(sub_655_2_n_85 | ~sub_655_2_n_67);
 assign sub_655_2_n_15 = ~(n_1506 | ~n_1479);
 assign sub_655_2_n_14 = ~(in1_65_15_ | ~n_1549);
 assign sub_655_2_n_13 = ~(in1_65_20_ | ~n_1593);
 assign sub_655_2_n_12 = ~(n_1476 | ~n_1579);
 assign sub_655_2_n_11 = ~(n_1535 & ~n_1515);
 assign sub_655_2_n_10 = ~(n_1513 | ~n_1555);
 assign sub_655_2_n_9 = (n_1514 & sub_655_2_n_60);
 assign sub_655_2_n_8 = ~(in1_65_19_ | ~n_1565);
 assign sub_655_2_n_7 = ~(n_1481 | ~n_1595);
 assign sub_655_2_n_6 = (n_1505 & sub_655_2_n_62);
 assign sub_655_2_n_5 = ~(in1_65_21_ | ~n_1591);
 assign sub_655_2_n_4 = ~(in1_65_17_ | ~n_1472);
 assign sub_655_2_n_3 = ~(n_1504 | ~n_1551);
 assign sub_655_2_n_2 = ~(n_1508 | ~n_1567);
 assign sub_655_2_n_1 = ~(n_1516 | ~n_1577);
 assign in1_67_1_ = (sub_655_2_n_54 ^ (n_1586 ^ n_1545));
 assign sub_676_2_n_188 = ~(sub_676_2_n_87 & (sub_676_2_n_185 | sub_676_2_n_11));
 assign in1_70_21_ = ~(sub_676_2_n_184 ^ sub_676_2_n_117);
 assign in1_70_19_ = (sub_676_2_n_183 ^ sub_676_2_n_23);
 assign sub_676_2_n_185 = ~(sub_676_2_n_38 | sub_676_2_n_140);
 assign sub_676_2_n_184 = ~(sub_676_2_n_95 & (sub_676_2_n_53 | sub_676_2_n_10));
 assign sub_676_2_n_183 = ~(sub_676_2_n_92 | (sub_676_2_n_178 & sub_676_2_n_86));
 assign in1_70_17_ = (sub_676_2_n_177 ^ sub_676_2_n_33);
 assign sub_676_2_n_181 = ~(sub_676_2_n_75 & (sub_676_2_n_175 | sub_676_2_n_89));
 assign in1_70_14_ = ~(sub_676_2_n_175 ^ sub_676_2_n_115);
 assign in1_70_24_ = ~(sub_676_2_n_50 | sub_676_2_n_158);
 assign sub_676_2_n_178 = ~(sub_676_2_n_141 & (sub_676_2_n_55 | sub_676_2_n_17));
 assign sub_676_2_n_177 = ~(sub_676_2_n_72 | (sub_676_2_n_56 & sub_676_2_n_0));
 assign sub_676_2_n_176 = ~(sub_676_2_n_172 & sub_676_2_n_137);
 assign sub_676_2_n_175 = ~(sub_676_2_n_131 | (sub_676_2_n_170 & sub_676_2_n_123));
 assign sub_676_2_n_174 = ~(sub_676_2_n_90 & (sub_676_2_n_171 | sub_676_2_n_2));
 assign sub_676_2_n_173 = ~(sub_676_2_n_99 & (sub_676_2_n_169 | sub_676_2_n_3));
 assign sub_676_2_n_172 = ~(sub_676_2_n_156 & (sub_676_2_n_166 | sub_676_2_n_138));
 assign sub_676_2_n_171 = ~sub_676_2_n_170;
 assign sub_676_2_n_170 = ~(sub_676_2_n_166 & sub_676_2_n_150);
 assign sub_676_2_n_169 = ~(sub_676_2_n_133 | (sub_676_2_n_162 & sub_676_2_n_107));
 assign sub_676_2_n_168 = ~(sub_676_2_n_94 & (sub_676_2_n_163 | sub_676_2_n_5));
 assign in1_70_8_ = ~(sub_676_2_n_163 ^ sub_676_2_n_29);
 assign sub_676_2_n_166 = ~(sub_676_2_n_162 & sub_676_2_n_136);
 assign sub_676_2_n_165 = ~(sub_676_2_n_77 & (sub_676_2_n_49 | sub_676_2_n_73));
 assign in1_70_5_ = (sub_676_2_n_161 ^ sub_676_2_n_116);
 assign sub_676_2_n_163 = ~sub_676_2_n_162;
 assign sub_676_2_n_162 = ~(sub_676_2_n_147 & (sub_676_2_n_159 | (sub_676_2_n_15 | sub_676_2_n_19)));
 assign sub_676_2_n_161 = ~(sub_676_2_n_98 & (sub_676_2_n_159 | sub_676_2_n_78));
 assign sub_676_2_n_160 = ~(sub_676_2_n_60 & (sub_676_2_n_153 | sub_676_2_n_7));
 assign sub_676_2_n_159 = ~(sub_676_2_n_157 | sub_676_2_n_128);
 assign sub_676_2_n_158 = ~(sub_676_2_n_154 & sub_676_2_n_149);
 assign sub_676_2_n_157 = ~(sub_676_2_n_153 | sub_676_2_n_28);
 assign sub_676_2_n_156 = ~(sub_676_2_n_146 | sub_676_2_n_155);
 assign sub_676_2_n_155 = ~(sub_676_2_n_150 | sub_676_2_n_138);
 assign sub_676_2_n_154 = ~(sub_676_2_n_148 & sub_676_2_n_139);
 assign sub_676_2_n_153 = ~(sub_676_2_n_152 | sub_676_2_n_6);
 assign sub_676_2_n_152 = ~(sub_676_2_n_145 & sub_676_2_n_51);
 assign in1_70_1_ = ~(in1_68_0_ ^ (n_1586 ^ sub_676_2_n_85));
 assign sub_676_2_n_150 = ~(sub_676_2_n_144 | sub_676_2_n_127);
 assign sub_676_2_n_149 = ~(sub_676_2_n_143 | sub_676_2_n_135);
 assign sub_676_2_n_148 = ~(sub_676_2_n_125 & (sub_676_2_n_141 | sub_676_2_n_122));
 assign sub_676_2_n_147 = ~(sub_676_2_n_142 | sub_676_2_n_129);
 assign sub_676_2_n_146 = ~(sub_676_2_n_126 & (sub_676_2_n_130 | sub_676_2_n_109));
 assign sub_676_2_n_145 = ~(sub_676_2_n_85 & ~n_1586);
 assign sub_676_2_n_144 = ~(sub_676_2_n_132 | sub_676_2_n_121);
 assign sub_676_2_n_143 = ~(sub_676_2_n_26 | ~sub_676_2_n_140);
 assign sub_676_2_n_142 = ~(sub_676_2_n_134 | sub_676_2_n_19);
 assign sub_676_2_n_137 = ~(sub_676_2_n_17 | sub_676_2_n_122);
 assign sub_676_2_n_136 = (sub_676_2_n_107 & sub_676_2_n_120);
 assign sub_676_2_n_135 = ~(sub_676_2_n_81 & (sub_676_2_n_87 | sub_676_2_n_12));
 assign sub_676_2_n_141 = ~(sub_676_2_n_103 | ~(sub_676_2_n_71 | sub_676_2_n_76));
 assign sub_676_2_n_140 = ~(sub_676_2_n_83 & (sub_676_2_n_95 | sub_676_2_n_8));
 assign sub_676_2_n_139 = ~(sub_676_2_n_26 | ~sub_676_2_n_112);
 assign sub_676_2_n_138 = ~(sub_676_2_n_123 & sub_676_2_n_108);
 assign sub_676_2_n_133 = ~sub_676_2_n_132;
 assign sub_676_2_n_131 = ~sub_676_2_n_130;
 assign sub_676_2_n_129 = ~(sub_676_2_n_80 & (sub_676_2_n_77 | sub_676_2_n_13));
 assign sub_676_2_n_128 = ~(sub_676_2_n_79 & (sub_676_2_n_60 | sub_676_2_n_93));
 assign sub_676_2_n_127 = ~(sub_676_2_n_84 & (sub_676_2_n_99 | sub_676_2_n_9));
 assign sub_676_2_n_126 = ~(sub_676_2_n_105 | sub_676_2_n_102);
 assign sub_676_2_n_125 = ~(sub_676_2_n_119 | sub_676_2_n_82);
 assign sub_676_2_n_134 = ~(sub_676_2_n_118 | sub_676_2_n_1);
 assign sub_676_2_n_132 = ~(sub_676_2_n_106 | sub_676_2_n_14);
 assign sub_676_2_n_130 = ~(sub_676_2_n_101 | ~(sub_676_2_n_90 | sub_676_2_n_91));
 assign sub_676_2_n_121 = ~sub_676_2_n_120;
 assign sub_676_2_n_119 = ~(sub_676_2_n_96 | ~sub_676_2_n_92);
 assign sub_676_2_n_118 = ~(sub_676_2_n_98 | sub_676_2_n_59);
 assign sub_676_2_n_117 = ~(sub_676_2_n_83 & ~sub_676_2_n_8);
 assign sub_676_2_n_124 = ~(sub_676_2_n_12 | ~sub_676_2_n_81);
 assign sub_676_2_n_123 = ~(sub_676_2_n_2 | sub_676_2_n_91);
 assign sub_676_2_n_116 = ~(sub_676_2_n_1 | sub_676_2_n_59);
 assign sub_676_2_n_122 = ~(sub_676_2_n_86 & sub_676_2_n_97);
 assign sub_676_2_n_120 = ~(sub_676_2_n_3 | sub_676_2_n_9);
 assign sub_676_2_n_115 = ~(sub_676_2_n_74 | sub_676_2_n_89);
 assign sub_676_2_n_109 = ~sub_676_2_n_108;
 assign sub_676_2_n_106 = ~(sub_676_2_n_94 | sub_676_2_n_88);
 assign sub_676_2_n_105 = ~(sub_676_2_n_100 | ~sub_676_2_n_74);
 assign in1_70_0_ = ~(sub_676_2_n_85 & ~(sub_676_2_n_61 & n_1599));
 assign sub_676_2_n_114 = ~(sub_676_2_n_14 | sub_676_2_n_88);
 assign sub_676_2_n_113 = ~(sub_676_2_n_102 | sub_676_2_n_100);
 assign sub_676_2_n_112 = ~(sub_676_2_n_10 | sub_676_2_n_8);
 assign sub_676_2_n_111 = ~(sub_676_2_n_101 | sub_676_2_n_91);
 assign sub_676_2_n_110 = ~(sub_676_2_n_9 | ~sub_676_2_n_84);
 assign sub_676_2_n_108 = ~(sub_676_2_n_89 | sub_676_2_n_100);
 assign sub_676_2_n_107 = ~(sub_676_2_n_5 | sub_676_2_n_88);
 assign sub_676_2_n_97 = ~sub_676_2_n_96;
 assign sub_676_2_n_103 = (sub_676_2_n_70 & in1_68_16_);
 assign sub_676_2_n_102 = (sub_676_2_n_66 & in1_68_14_);
 assign sub_676_2_n_101 = (sub_676_2_n_62 & in1_68_12_);
 assign sub_676_2_n_100 = ~(in1_68_14_ | sub_676_2_n_66);
 assign sub_676_2_n_99 = ~(in1_68_9_ & ~n_1551);
 assign sub_676_2_n_98 = ~(in1_68_3_ & ~n_1535);
 assign sub_676_2_n_96 = ~(in1_68_18_ | sub_676_2_n_64);
 assign sub_676_2_n_95 = ~(in1_68_19_ & ~n_1565);
 assign sub_676_2_n_94 = ~(in1_68_7_ & ~n_1479);
 assign sub_676_2_n_93 = ~(in1_68_2_ | sub_676_2_n_68);
 assign sub_676_2_n_92 = (sub_676_2_n_65 & in1_68_17_);
 assign sub_676_2_n_91 = ~(in1_68_12_ | sub_676_2_n_62);
 assign sub_676_2_n_90 = ~(in1_68_11_ & ~n_1595);
 assign sub_676_2_n_89 = ~(sub_676_2_n_58 | sub_676_2_n_67);
 assign sub_676_2_n_88 = ~(in1_68_8_ | sub_676_2_n_63);
 assign sub_676_2_n_87 = ~(in1_68_21_ & ~n_1591);
 assign sub_676_2_n_86 = (in1_68_17_ | sub_676_2_n_65);
 assign sub_676_2_n_85 = ~(n_1543 & ~n_1599);
 assign sub_676_2_n_78 = ~sub_676_2_n_4;
 assign sub_676_2_n_75 = ~sub_676_2_n_74;
 assign sub_676_2_n_72 = ~sub_676_2_n_71;
 assign sub_676_2_n_84 = ~(in1_68_10_ & ~n_1555);
 assign sub_676_2_n_83 = ~(in1_68_20_ & ~n_1593);
 assign sub_676_2_n_82 = (sub_676_2_n_64 & in1_68_18_);
 assign sub_676_2_n_81 = ~(in1_68_22_ & ~n_1403);
 assign sub_676_2_n_80 = ~(in1_68_6_ & ~n_1527);
 assign sub_676_2_n_79 = ~(in1_68_2_ & ~n_1579);
 assign sub_676_2_n_60 = ~(in1_68_1_ & ~n_1477);
 assign sub_676_2_n_77 = ~(in1_68_5_ & ~n_1567);
 assign sub_676_2_n_76 = ~(in1_68_16_ | sub_676_2_n_70);
 assign sub_676_2_n_74 = (sub_676_2_n_67 & in1_68_13_);
 assign sub_676_2_n_59 = ~(in1_68_4_ | sub_676_2_n_69);
 assign sub_676_2_n_73 = ~(in1_68_5_ | ~n_1567);
 assign sub_676_2_n_71 = ~(in1_68_15_ & ~n_1549);
 assign sub_676_2_n_70 = ~n_1562;
 assign sub_676_2_n_69 = ~n_1569;
 assign sub_676_2_n_68 = ~n_1579;
 assign sub_676_2_n_67 = ~n_1577;
 assign sub_676_2_n_66 = ~n_1495;
 assign sub_676_2_n_65 = ~n_1472;
 assign sub_676_2_n_64 = ~n_1558;
 assign sub_676_2_n_63 = ~n_1589;
 assign sub_676_2_n_62 = ~n_1581;
 assign sub_676_2_n_61 = ~n_1543;
 assign sub_676_2_n_58 = in1_68_13_;
 assign sub_676_2_n_57 = in1_68_7_;
 assign sub_676_2_n_56 = ~sub_676_2_n_55;
 assign sub_676_2_n_55 = ~sub_676_2_n_172;
 assign in1_70_18_ = ~(sub_676_2_n_178 ^ sub_676_2_n_27);
 assign sub_676_2_n_53 = ~(sub_676_2_n_148 | ~sub_676_2_n_176);
 assign in1_70_10_ = ~(sub_676_2_n_169 ^ sub_676_2_n_32);
 assign sub_676_2_n_51 = ~(in1_68_0_ & sub_676_2_n_85);
 assign sub_676_2_n_50 = ~(sub_676_2_n_176 | ~sub_676_2_n_139);
 assign sub_676_2_n_49 = (sub_676_2_n_134 & (sub_676_2_n_159 | sub_676_2_n_15));
 assign in1_70_23_ = (sub_676_2_n_188 ^ sub_676_2_n_124);
 assign in1_70_4_ = ~(sub_676_2_n_159 ^ sub_676_2_n_31);
 assign in1_70_22_ = ~(sub_676_2_n_185 ^ sub_676_2_n_24);
 assign in1_70_2_ = ~(sub_676_2_n_153 ^ sub_676_2_n_20);
 assign in1_70_6_ = ~(sub_676_2_n_49 ^ sub_676_2_n_18);
 assign in1_70_20_ = ~(sub_676_2_n_53 ^ sub_676_2_n_30);
 assign in1_70_9_ = (sub_676_2_n_168 ^ sub_676_2_n_114);
 assign in1_70_16_ = (sub_676_2_n_56 ^ sub_676_2_n_16);
 assign in1_70_3_ = (sub_676_2_n_160 ^ sub_676_2_n_21);
 assign in1_70_15_ = (sub_676_2_n_181 ^ sub_676_2_n_113);
 assign sub_676_2_n_38 = ~(sub_676_2_n_53 | ~sub_676_2_n_112);
 assign in1_70_13_ = (sub_676_2_n_174 ^ sub_676_2_n_111);
 assign in1_70_11_ = (sub_676_2_n_173 ^ sub_676_2_n_110);
 assign in1_70_12_ = (sub_676_2_n_170 ^ sub_676_2_n_25);
 assign in1_70_7_ = (sub_676_2_n_165 ^ sub_676_2_n_22);
 assign sub_676_2_n_33 = (sub_676_2_n_103 | sub_676_2_n_76);
 assign sub_676_2_n_32 = ~(sub_676_2_n_3 | ~sub_676_2_n_99);
 assign sub_676_2_n_31 = ~(sub_676_2_n_78 | ~sub_676_2_n_98);
 assign sub_676_2_n_30 = ~(sub_676_2_n_10 | ~sub_676_2_n_95);
 assign sub_676_2_n_29 = ~(sub_676_2_n_5 | ~sub_676_2_n_94);
 assign sub_676_2_n_28 = (sub_676_2_n_93 | sub_676_2_n_7);
 assign sub_676_2_n_27 = ~(sub_676_2_n_86 & ~sub_676_2_n_92);
 assign sub_676_2_n_26 = (sub_676_2_n_12 | sub_676_2_n_11);
 assign sub_676_2_n_25 = ~(sub_676_2_n_2 | ~sub_676_2_n_90);
 assign sub_676_2_n_24 = ~(sub_676_2_n_11 | ~sub_676_2_n_87);
 assign sub_676_2_n_23 = ~(sub_676_2_n_97 & ~sub_676_2_n_82);
 assign sub_676_2_n_22 = ~(sub_676_2_n_13 | ~sub_676_2_n_80);
 assign sub_676_2_n_21 = ~(sub_676_2_n_93 | ~sub_676_2_n_79);
 assign sub_676_2_n_20 = ~(sub_676_2_n_7 | ~sub_676_2_n_60);
 assign sub_676_2_n_19 = (sub_676_2_n_13 | sub_676_2_n_73);
 assign sub_676_2_n_18 = ~(sub_676_2_n_73 | ~sub_676_2_n_77);
 assign sub_676_2_n_17 = ~(sub_676_2_n_0 & ~sub_676_2_n_76);
 assign sub_676_2_n_16 = ~(sub_676_2_n_72 | ~sub_676_2_n_0);
 assign sub_676_2_n_15 = ~(sub_676_2_n_4 & ~sub_676_2_n_59);
 assign sub_676_2_n_14 = (in1_68_8_ & sub_676_2_n_63);
 assign sub_676_2_n_13 = ~(in1_68_6_ | ~n_1527);
 assign sub_676_2_n_12 = ~(in1_68_22_ | ~n_1403);
 assign sub_676_2_n_11 = ~(in1_68_21_ | ~n_1591);
 assign sub_676_2_n_10 = ~(in1_68_19_ | ~n_1565);
 assign sub_676_2_n_9 = ~(in1_68_10_ | ~n_1555);
 assign sub_676_2_n_8 = ~(in1_68_20_ | ~n_1593);
 assign sub_676_2_n_7 = ~(in1_68_1_ | ~n_1477);
 assign sub_676_2_n_6 = ~(n_1586 | ~in1_68_0_);
 assign sub_676_2_n_5 = ~(sub_676_2_n_57 | ~n_1479);
 assign sub_676_2_n_4 = ~(n_1535 & ~in1_68_3_);
 assign sub_676_2_n_3 = ~(in1_68_9_ | ~n_1551);
 assign sub_676_2_n_2 = ~(in1_68_11_ | ~n_1595);
 assign sub_676_2_n_1 = (in1_68_4_ & sub_676_2_n_69);
 assign sub_676_2_n_0 = ~(n_1549 & ~in1_68_15_);
 assign sub_697_2_n_206 = ~(sub_697_2_n_203 | sub_697_2_n_71);
 assign in1_73_21_ = (sub_697_2_n_200 ^ sub_697_2_n_120);
 assign in1_73_19_ = (sub_697_2_n_17 ^ sub_697_2_n_119);
 assign sub_697_2_n_203 = ~(sub_697_2_n_201 | sub_697_2_n_64);
 assign sub_697_2_n_202 = ~(sub_697_2_n_189 | in1_71_23_);
 assign sub_697_2_n_201 = ~(sub_697_2_n_196 | sub_697_2_n_143);
 assign sub_697_2_n_200 = ~(sub_697_2_n_195 | sub_697_2_n_94);
 assign in1_73_20_ = ~(sub_697_2_n_193 & ~sub_697_2_n_194);
 assign in1_73_17_ = (sub_697_2_n_187 ^ sub_697_2_n_21);
 assign in1_73_18_ = (sub_697_2_n_40 ^ sub_697_2_n_118);
 assign sub_697_2_n_196 = ~(sub_697_2_n_45 | sub_697_2_n_111);
 assign sub_697_2_n_195 = ~(sub_697_2_n_45 | sub_697_2_n_6);
 assign sub_697_2_n_194 = ~(sub_697_2_n_45 | sub_697_2_n_127);
 assign sub_697_2_n_193 = ~(sub_697_2_n_45 & sub_697_2_n_127);
 assign sub_697_2_n_192 = ~(sub_697_2_n_40 | sub_697_2_n_83);
 assign sub_697_2_n_191 = ~(sub_697_2_n_188 | sub_697_2_n_91);
 assign in1_73_14_ = ~(sub_697_2_n_42 ^ sub_697_2_n_103);
 assign sub_697_2_n_189 = ~(sub_697_2_n_163 & (sub_697_2_n_185 | sub_697_2_n_145));
 assign sub_697_2_n_188 = ~(sub_697_2_n_42 | sub_697_2_n_2);
 assign sub_697_2_n_187 = ~(sub_697_2_n_96 | ~(sub_697_2_n_180 | sub_697_2_n_65));
 assign in1_73_16_ = (sub_697_2_n_180 ^ sub_697_2_n_102);
 assign sub_697_2_n_185 = ~(sub_697_2_n_179 & sub_697_2_n_36);
 assign sub_697_2_n_184 = ~(sub_697_2_n_182 | sub_697_2_n_62);
 assign sub_697_2_n_183 = ~(sub_697_2_n_181 | sub_697_2_n_89);
 assign sub_697_2_n_182 = ~(sub_697_2_n_43 | sub_697_2_n_7);
 assign sub_697_2_n_181 = ~(sub_697_2_n_41 | sub_697_2_n_5);
 assign sub_697_2_n_180 = ~sub_697_2_n_179;
 assign sub_697_2_n_179 = ~(sub_697_2_n_162 & (sub_697_2_n_173 | (sub_697_2_n_32 | sub_697_2_n_142)));
 assign sub_697_2_n_178 = ~(sub_697_2_n_87 | ~(sub_697_2_n_173 | sub_697_2_n_79));
 assign in1_73_8_ = ~(sub_697_2_n_173 ^ sub_697_2_n_104);
 assign sub_697_2_n_176 = ~(sub_697_2_n_173 | sub_697_2_n_32);
 assign sub_697_2_n_175 = ~(sub_697_2_n_69 | (sub_697_2_n_171 & sub_697_2_n_9));
 assign in1_73_6_ = (sub_697_2_n_171 ^ sub_697_2_n_19);
 assign sub_697_2_n_173 = ~(sub_697_2_n_172 | sub_697_2_n_153);
 assign sub_697_2_n_172 = ~(sub_697_2_n_167 | (sub_697_2_n_16 | sub_697_2_n_13));
 assign sub_697_2_n_171 = ~(sub_697_2_n_140 & (sub_697_2_n_167 | sub_697_2_n_16));
 assign sub_697_2_n_170 = ~(sub_697_2_n_81 | (sub_697_2_n_168 & sub_697_2_n_1));
 assign in1_73_2_ = ~(sub_697_2_n_166 & ~sub_697_2_n_165);
 assign sub_697_2_n_168 = ~sub_697_2_n_167;
 assign sub_697_2_n_167 = ~(sub_697_2_n_164 | sub_697_2_n_141);
 assign sub_697_2_n_166 = ~(sub_697_2_n_159 & sub_697_2_n_126);
 assign sub_697_2_n_165 = ~(sub_697_2_n_159 | sub_697_2_n_126);
 assign sub_697_2_n_164 = ~(sub_697_2_n_159 | sub_697_2_n_14);
 assign sub_697_2_n_163 = ~(sub_697_2_n_160 | sub_697_2_n_154);
 assign sub_697_2_n_162 = ~(sub_697_2_n_161 | sub_697_2_n_152);
 assign sub_697_2_n_161 = ~(sub_697_2_n_155 | sub_697_2_n_142);
 assign sub_697_2_n_160 = ~(sub_697_2_n_156 | sub_697_2_n_145);
 assign sub_697_2_n_159 = ~(sub_697_2_n_158 | sub_697_2_n_77);
 assign sub_697_2_n_158 = ~(sub_697_2_n_150 & sub_697_2_n_151);
 assign in1_73_1_ = ~((sub_697_2_n_146 & ~sub_697_2_n_101) | (sub_697_2_n_60 & sub_697_2_n_101));
 assign sub_697_2_n_156 = ~(sub_697_2_n_148 | sub_697_2_n_136);
 assign sub_697_2_n_155 = ~(sub_697_2_n_147 | sub_697_2_n_135);
 assign sub_697_2_n_154 = ~(sub_697_2_n_149 & sub_697_2_n_133);
 assign sub_697_2_n_153 = ~(sub_697_2_n_134 & (sub_697_2_n_140 | sub_697_2_n_13));
 assign sub_697_2_n_152 = ~(sub_697_2_n_137 & (sub_697_2_n_144 | sub_697_2_n_125));
 assign sub_697_2_n_151 = ~(in1_71_0_ & ~sub_697_2_n_146);
 assign sub_697_2_n_150 = ~(sub_697_2_n_60 & ~n_1586);
 assign sub_697_2_n_149 = ~(sub_697_2_n_143 & sub_697_2_n_109);
 assign sub_697_2_n_148 = ~(sub_697_2_n_138 | sub_697_2_n_18);
 assign sub_697_2_n_147 = ~(sub_697_2_n_139 | sub_697_2_n_20);
 assign sub_697_2_n_146 = ~sub_697_2_n_60;
 assign sub_697_2_n_141 = ~(sub_697_2_n_100 & (sub_697_2_n_84 | sub_697_2_n_12));
 assign sub_697_2_n_145 = ~(sub_697_2_n_109 & ~sub_697_2_n_111);
 assign sub_697_2_n_144 = ~(sub_697_2_n_122 | sub_697_2_n_97);
 assign sub_697_2_n_143 = ~(sub_697_2_n_76 & (sub_697_2_n_93 | sub_697_2_n_8));
 assign sub_697_2_n_142 = ~(sub_697_2_n_129 & sub_697_2_n_124);
 assign sub_697_2_n_137 = ~(sub_697_2_n_75 | ~(sub_697_2_n_90 | sub_697_2_n_92));
 assign sub_697_2_n_136 = ~(sub_697_2_n_99 & (sub_697_2_n_82 | sub_697_2_n_3));
 assign sub_697_2_n_135 = ~(sub_697_2_n_74 & (sub_697_2_n_88 | sub_697_2_n_0));
 assign sub_697_2_n_134 = ~(sub_697_2_n_73 | ~(sub_697_2_n_68 | sub_697_2_n_48));
 assign sub_697_2_n_133 = ~(sub_697_2_n_123 | sub_697_2_n_11);
 assign sub_697_2_n_140 = ~(sub_697_2_n_121 | sub_697_2_n_72);
 assign sub_697_2_n_139 = ~(sub_697_2_n_107 | sub_697_2_n_10);
 assign sub_697_2_n_138 = ~(sub_697_2_n_106 | sub_697_2_n_98);
 assign sub_697_2_n_125 = ~sub_697_2_n_124;
 assign sub_697_2_n_123 = ~(sub_697_2_n_4 | ~sub_697_2_n_71);
 assign sub_697_2_n_122 = ~(sub_697_2_n_61 | sub_697_2_n_66);
 assign sub_697_2_n_121 = ~(sub_697_2_n_80 | sub_697_2_n_49);
 assign sub_697_2_n_132 = ~(sub_697_2_n_73 | sub_697_2_n_48);
 assign sub_697_2_n_131 = ~(sub_697_2_n_72 | sub_697_2_n_49);
 assign sub_697_2_n_130 = ~(sub_697_2_n_11 | sub_697_2_n_4);
 assign sub_697_2_n_129 = ~(sub_697_2_n_7 | sub_697_2_n_66);
 assign sub_697_2_n_128 = ~(sub_697_2_n_71 | sub_697_2_n_64);
 assign sub_697_2_n_120 = ~(sub_697_2_n_76 & ~sub_697_2_n_8);
 assign sub_697_2_n_127 = ~(sub_697_2_n_94 | sub_697_2_n_6);
 assign sub_697_2_n_126 = ~(sub_697_2_n_85 | sub_697_2_n_63);
 assign sub_697_2_n_119 = ~(sub_697_2_n_99 & ~sub_697_2_n_3);
 assign sub_697_2_n_118 = ~(sub_697_2_n_82 & ~sub_697_2_n_83);
 assign sub_697_2_n_124 = ~(sub_697_2_n_2 | sub_697_2_n_92);
 assign sub_697_2_n_107 = ~(sub_697_2_n_86 | sub_697_2_n_67);
 assign sub_697_2_n_106 = ~(sub_697_2_n_95 | sub_697_2_n_70);
 assign in1_73_0_ = ~(sub_697_2_n_60 & ~(sub_697_2_n_54 & n_1572));
 assign sub_697_2_n_117 = ~(sub_697_2_n_89 | sub_697_2_n_5);
 assign sub_697_2_n_104 = ~(sub_697_2_n_87 | sub_697_2_n_79);
 assign sub_697_2_n_103 = ~(sub_697_2_n_91 | sub_697_2_n_2);
 assign sub_697_2_n_116 = ~(sub_697_2_n_79 | sub_697_2_n_67);
 assign sub_697_2_n_115 = ~(sub_697_2_n_10 | sub_697_2_n_67);
 assign sub_697_2_n_114 = ~(sub_697_2_n_0 | ~sub_697_2_n_74);
 assign sub_697_2_n_113 = ~(sub_697_2_n_62 | sub_697_2_n_7);
 assign sub_697_2_n_102 = (sub_697_2_n_96 | sub_697_2_n_65);
 assign sub_697_2_n_112 = ~(sub_697_2_n_65 | sub_697_2_n_70);
 assign sub_697_2_n_111 = (sub_697_2_n_6 | sub_697_2_n_8);
 assign sub_697_2_n_110 = ~(sub_697_2_n_97 | sub_697_2_n_66);
 assign sub_697_2_n_109 = ~(sub_697_2_n_64 | sub_697_2_n_4);
 assign sub_697_2_n_108 = ~(sub_697_2_n_75 | sub_697_2_n_92);
 assign sub_697_2_n_101 = ~(sub_697_2_n_77 | sub_697_2_n_78);
 assign sub_697_2_n_96 = ~sub_697_2_n_95;
 assign sub_697_2_n_94 = ~sub_697_2_n_93;
 assign sub_697_2_n_91 = ~sub_697_2_n_90;
 assign sub_697_2_n_89 = ~sub_697_2_n_88;
 assign sub_697_2_n_87 = ~sub_697_2_n_86;
 assign sub_697_2_n_85 = ~sub_697_2_n_84;
 assign sub_697_2_n_81 = ~sub_697_2_n_80;
 assign sub_697_2_n_78 = ~(in1_71_0_ | ~n_1586);
 assign sub_697_2_n_100 = ~(in1_71_2_ & ~n_1579);
 assign sub_697_2_n_99 = ~(in1_71_18_ & ~n_1558);
 assign sub_697_2_n_98 = (sub_697_2_n_51 & in1_71_16_);
 assign sub_697_2_n_97 = (sub_697_2_n_53 & in1_71_12_);
 assign sub_697_2_n_95 = ~(in1_71_15_ & ~n_1549);
 assign sub_697_2_n_93 = ~(in1_71_19_ & ~n_1565);
 assign sub_697_2_n_92 = ~(in1_71_14_ | sub_697_2_n_52);
 assign sub_697_2_n_90 = ~(in1_71_13_ & ~n_1577);
 assign sub_697_2_n_88 = ~(in1_71_9_ & ~n_1551);
 assign sub_697_2_n_86 = ~(in1_71_7_ & ~n_1479);
 assign sub_697_2_n_84 = ~(in1_71_1_ & ~n_1477);
 assign sub_697_2_n_83 = ~(in1_71_17_ | ~n_1472);
 assign sub_697_2_n_82 = ~(in1_71_17_ & ~n_1472);
 assign sub_697_2_n_80 = ~(in1_71_3_ & ~n_1535);
 assign sub_697_2_n_79 = ~(in1_71_7_ | ~n_1479);
 assign sub_697_2_n_69 = ~sub_697_2_n_68;
 assign sub_697_2_n_62 = ~sub_697_2_n_61;
 assign sub_697_2_n_77 = ~(sub_697_2_n_55 | ~sub_697_2_n_56);
 assign sub_697_2_n_76 = ~(in1_71_20_ & ~n_1593);
 assign sub_697_2_n_75 = (sub_697_2_n_52 & in1_71_14_);
 assign sub_697_2_n_74 = ~(in1_71_10_ & ~n_1555);
 assign sub_697_2_n_73 = (sub_697_2_n_57 & in1_71_6_);
 assign sub_697_2_n_72 = (sub_697_2_n_58 & in1_71_4_);
 assign sub_697_2_n_49 = ~(in1_71_4_ | sub_697_2_n_58);
 assign sub_697_2_n_71 = (sub_697_2_n_50 & in1_71_21_);
 assign sub_697_2_n_70 = ~(in1_71_16_ | sub_697_2_n_51);
 assign sub_697_2_n_68 = ~(in1_71_5_ & ~n_1567);
 assign sub_697_2_n_67 = ~(in1_71_8_ | sub_697_2_n_59);
 assign sub_697_2_n_66 = ~(in1_71_12_ | sub_697_2_n_53);
 assign sub_697_2_n_65 = ~(in1_71_15_ | ~n_1549);
 assign sub_697_2_n_64 = ~(in1_71_21_ | sub_697_2_n_50);
 assign sub_697_2_n_63 = ~(in1_71_1_ | ~n_1477);
 assign sub_697_2_n_61 = ~(in1_71_11_ & ~n_1595);
 assign sub_697_2_n_48 = ~(in1_71_6_ | sub_697_2_n_57);
 assign sub_697_2_n_60 = ~(n_1543 & ~n_1572);
 assign sub_697_2_n_59 = ~n_1589;
 assign sub_697_2_n_58 = ~n_1569;
 assign sub_697_2_n_57 = ~n_1527;
 assign sub_697_2_n_56 = ~n_1586;
 assign sub_697_2_n_55 = ~in1_71_0_;
 assign sub_697_2_n_54 = ~n_1543;
 assign sub_697_2_n_53 = ~n_1581;
 assign sub_697_2_n_52 = ~n_1495;
 assign sub_697_2_n_51 = ~n_1562;
 assign sub_697_2_n_50 = ~n_1591;
 assign in1_73_24_ = (sub_697_2_n_202 | sub_697_2_n_46);
 assign sub_697_2_n_46 = (sub_697_2_n_189 & in1_71_23_);
 assign sub_697_2_n_45 = (sub_697_2_n_185 & sub_697_2_n_156);
 assign sub_697_2_n_44 = ~(sub_697_2_n_85 | ~(sub_697_2_n_159 | sub_697_2_n_63));
 assign sub_697_2_n_43 = ~(sub_697_2_n_176 | ~sub_697_2_n_155);
 assign sub_697_2_n_42 = ~(sub_697_2_n_35 | ~sub_697_2_n_144);
 assign sub_697_2_n_41 = ~(sub_697_2_n_29 | ~sub_697_2_n_139);
 assign sub_697_2_n_40 = ~(sub_697_2_n_25 | ~sub_697_2_n_138);
 assign in1_73_7_ = ~(sub_697_2_n_175 ^ sub_697_2_n_132);
 assign in1_73_5_ = ~(sub_697_2_n_170 ^ sub_697_2_n_131);
 assign in1_73_23_ = ~(sub_697_2_n_206 ^ sub_697_2_n_130);
 assign sub_697_2_n_36 = ~(sub_697_2_n_18 | ~sub_697_2_n_112);
 assign sub_697_2_n_35 = ~(sub_697_2_n_43 | ~sub_697_2_n_129);
 assign in1_73_3_ = ~(sub_697_2_n_44 ^ sub_697_2_n_22);
 assign in1_73_22_ = ~(sub_697_2_n_201 ^ sub_697_2_n_128);
 assign sub_697_2_n_32 = ~(sub_697_2_n_116 & ~sub_697_2_n_20);
 assign in1_73_4_ = ~(sub_697_2_n_167 ^ sub_697_2_n_15);
 assign in1_73_10_ = ~(sub_697_2_n_41 ^ sub_697_2_n_117);
 assign sub_697_2_n_29 = ~(sub_697_2_n_173 | ~sub_697_2_n_116);
 assign in1_73_9_ = ~(sub_697_2_n_178 ^ sub_697_2_n_115);
 assign in1_73_11_ = ~(sub_697_2_n_183 ^ sub_697_2_n_114);
 assign in1_73_12_ = ~(sub_697_2_n_43 ^ sub_697_2_n_113);
 assign sub_697_2_n_25 = ~(sub_697_2_n_180 | ~sub_697_2_n_112);
 assign in1_73_13_ = ~(sub_697_2_n_184 ^ sub_697_2_n_110);
 assign in1_73_15_ = ~(sub_697_2_n_191 ^ sub_697_2_n_108);
 assign sub_697_2_n_22 = ~(sub_697_2_n_12 | ~sub_697_2_n_100);
 assign sub_697_2_n_21 = (sub_697_2_n_98 | sub_697_2_n_70);
 assign sub_697_2_n_20 = (sub_697_2_n_0 | sub_697_2_n_5);
 assign sub_697_2_n_19 = ~(sub_697_2_n_69 | ~sub_697_2_n_9);
 assign sub_697_2_n_18 = (sub_697_2_n_3 | sub_697_2_n_83);
 assign sub_697_2_n_17 = ~(sub_697_2_n_192 | ~sub_697_2_n_82);
 assign sub_697_2_n_16 = ~(sub_697_2_n_1 & ~sub_697_2_n_49);
 assign sub_697_2_n_15 = ~(sub_697_2_n_81 | ~sub_697_2_n_1);
 assign sub_697_2_n_14 = (sub_697_2_n_12 | sub_697_2_n_63);
 assign sub_697_2_n_13 = ~(sub_697_2_n_9 & ~sub_697_2_n_48);
 assign sub_697_2_n_12 = ~(in1_71_2_ | ~n_1579);
 assign sub_697_2_n_11 = ~(n_1403 | ~in1_71_22_);
 assign sub_697_2_n_10 = (in1_71_8_ & sub_697_2_n_59);
 assign sub_697_2_n_9 = ~(n_1567 & ~in1_71_5_);
 assign sub_697_2_n_8 = ~(in1_71_20_ | ~n_1593);
 assign sub_697_2_n_7 = ~(in1_71_11_ | ~n_1595);
 assign sub_697_2_n_6 = ~(in1_71_19_ | ~n_1565);
 assign sub_697_2_n_5 = ~(in1_71_9_ | ~n_1551);
 assign sub_697_2_n_4 = ~(in1_71_22_ | ~n_1403);
 assign sub_697_2_n_3 = ~(in1_71_18_ | ~n_1558);
 assign sub_697_2_n_2 = ~(in1_71_13_ | ~n_1577);
 assign sub_697_2_n_1 = ~(n_1535 & ~in1_71_3_);
 assign sub_697_2_n_0 = ~(in1_71_10_ | ~n_1555);
 assign sub_718_2_n_202 = ~(sub_718_2_n_73 | (sub_718_2_n_200 & sub_718_2_n_7));
 assign in1_76_19_ = (sub_718_2_n_198 ^ sub_718_2_n_106);
 assign sub_718_2_n_200 = ~(sub_718_2_n_138 & (sub_718_2_n_191 | sub_718_2_n_20));
 assign sub_718_2_n_199 = ~(sub_718_2_n_71 | (sub_718_2_n_192 & sub_718_2_n_3));
 assign sub_718_2_n_198 = ~(sub_718_2_n_79 & (sub_718_2_n_42 | sub_718_2_n_8));
 assign sub_718_2_n_197 = ~(sub_718_2_n_97 & (sub_718_2_n_193 | sub_718_2_n_6));
 assign in1_76_18_ = ~(sub_718_2_n_42 ^ sub_718_2_n_15);
 assign in1_76_17_ = ~(sub_718_2_n_189 ^ sub_718_2_n_107);
 assign in1_76_24_ = ~(sub_718_2_n_2 & sub_718_2_n_190);
 assign sub_718_2_n_192 = ~sub_718_2_n_191;
 assign sub_718_2_n_190 = ~(sub_718_2_n_183 & in1_74_23_);
 assign sub_718_2_n_189 = ~(sub_718_2_n_66 | (sub_718_2_n_181 & sub_718_2_n_4));
 assign sub_718_2_n_193 = ~(sub_718_2_n_140 | (sub_718_2_n_180 & sub_718_2_n_128));
 assign sub_718_2_n_191 = ~(sub_718_2_n_43 | sub_718_2_n_156);
 assign in1_76_12_ = ~(sub_718_2_n_180 ^ sub_718_2_n_104);
 assign in1_76_16_ = ~(sub_718_2_n_46 ^ sub_718_2_n_13);
 assign sub_718_2_n_186 = ~(sub_718_2_n_95 & (sub_718_2_n_179 | sub_718_2_n_5));
 assign sub_718_2_n_185 = ~(sub_718_2_n_92 & (sub_718_2_n_178 | sub_718_2_n_75));
 assign sub_718_2_n_184 = ~(sub_718_2_n_46 | sub_718_2_n_21);
 assign sub_718_2_n_183 = ~sub_718_2_n_182;
 assign sub_718_2_n_182 = ~(sub_718_2_n_168 | (sub_718_2_n_174 & sub_718_2_n_152));
 assign sub_718_2_n_181 = ~sub_718_2_n_46;
 assign sub_718_2_n_179 = ~sub_718_2_n_180;
 assign sub_718_2_n_180 = ~(sub_718_2_n_159 & (sub_718_2_n_173 | sub_718_2_n_148));
 assign sub_718_2_n_178 = ~(sub_718_2_n_136 | (sub_718_2_n_172 & sub_718_2_n_113));
 assign sub_718_2_n_177 = ~(sub_718_2_n_76 & (sub_718_2_n_173 | sub_718_2_n_10));
 assign in1_76_8_ = ~(sub_718_2_n_173 ^ sub_718_2_n_14);
 assign sub_718_2_n_175 = ~(sub_718_2_n_93 & (sub_718_2_n_170 | sub_718_2_n_96));
 assign sub_718_2_n_174 = ~(sub_718_2_n_173 | sub_718_2_n_44);
 assign sub_718_2_n_172 = ~sub_718_2_n_173;
 assign sub_718_2_n_173 = ~(sub_718_2_n_171 | sub_718_2_n_158);
 assign sub_718_2_n_171 = ~(sub_718_2_n_166 | (sub_718_2_n_130 | sub_718_2_n_19));
 assign sub_718_2_n_170 = ~(sub_718_2_n_142 | (sub_718_2_n_165 & sub_718_2_n_131));
 assign sub_718_2_n_169 = ~(sub_718_2_n_91 | (sub_718_2_n_165 & sub_718_2_n_9));
 assign sub_718_2_n_168 = ~(sub_718_2_n_162 & (sub_718_2_n_163 | sub_718_2_n_151));
 assign sub_718_2_n_167 = ~(sub_718_2_n_68 | (sub_718_2_n_161 & sub_718_2_n_0));
 assign sub_718_2_n_165 = ~sub_718_2_n_166;
 assign sub_718_2_n_166 = ~(sub_718_2_n_164 | sub_718_2_n_133);
 assign sub_718_2_n_164 = ~(sub_718_2_n_154 | sub_718_2_n_18);
 assign sub_718_2_n_163 = ~(sub_718_2_n_160 | sub_718_2_n_157);
 assign sub_718_2_n_162 = ~(sub_718_2_n_155 | (sub_718_2_n_156 & sub_718_2_n_147));
 assign sub_718_2_n_161 = ~sub_718_2_n_154;
 assign sub_718_2_n_160 = ~(sub_718_2_n_159 | sub_718_2_n_149);
 assign sub_718_2_n_159 = ~(sub_718_2_n_153 | sub_718_2_n_134);
 assign sub_718_2_n_158 = ~(sub_718_2_n_144 & (sub_718_2_n_141 | sub_718_2_n_19));
 assign sub_718_2_n_157 = ~(sub_718_2_n_145 & (sub_718_2_n_139 | sub_718_2_n_126));
 assign sub_718_2_n_156 = ~(sub_718_2_n_143 & (sub_718_2_n_137 | sub_718_2_n_12));
 assign sub_718_2_n_155 = ~(sub_718_2_n_132 & (sub_718_2_n_138 | sub_718_2_n_25));
 assign sub_718_2_n_154 = ~(sub_718_2_n_150 | sub_718_2_n_82);
 assign sub_718_2_n_153 = ~(sub_718_2_n_135 | sub_718_2_n_17);
 assign sub_718_2_n_152 = ~sub_718_2_n_151;
 assign sub_718_2_n_151 = ~(sub_718_2_n_146 & sub_718_2_n_147);
 assign sub_718_2_n_150 = ~(sub_718_2_n_87 | ~sub_718_2_n_64);
 assign sub_718_2_n_148 = ~sub_718_2_n_33;
 assign sub_718_2_n_145 = ~(sub_718_2_n_121 | sub_718_2_n_88);
 assign sub_718_2_n_144 = ~(sub_718_2_n_122 | sub_718_2_n_84);
 assign sub_718_2_n_143 = ~(sub_718_2_n_117 | sub_718_2_n_102);
 assign sub_718_2_n_149 = ~(sub_718_2_n_128 & sub_718_2_n_125);
 assign sub_718_2_n_147 = ~(sub_718_2_n_20 | sub_718_2_n_25);
 assign sub_718_2_n_146 = ~(sub_718_2_n_21 | sub_718_2_n_12);
 assign sub_718_2_n_142 = ~sub_718_2_n_141;
 assign sub_718_2_n_140 = ~sub_718_2_n_139;
 assign sub_718_2_n_136 = ~sub_718_2_n_135;
 assign sub_718_2_n_134 = ~(sub_718_2_n_101 & (sub_718_2_n_92 | sub_718_2_n_1));
 assign sub_718_2_n_133 = ~(sub_718_2_n_103 & (sub_718_2_n_67 | sub_718_2_n_81));
 assign sub_718_2_n_132 = ~(sub_718_2_n_85 | ~(sub_718_2_n_72 | sub_718_2_n_51));
 assign sub_718_2_n_141 = ~(sub_718_2_n_118 | sub_718_2_n_86);
 assign sub_718_2_n_139 = ~(sub_718_2_n_123 | sub_718_2_n_100);
 assign sub_718_2_n_138 = ~(sub_718_2_n_83 | ~(sub_718_2_n_70 | sub_718_2_n_50));
 assign sub_718_2_n_137 = ~(sub_718_2_n_120 | sub_718_2_n_98);
 assign sub_718_2_n_135 = ~(sub_718_2_n_119 | sub_718_2_n_99);
 assign sub_718_2_n_131 = ~sub_718_2_n_130;
 assign sub_718_2_n_126 = ~sub_718_2_n_125;
 assign sub_718_2_n_123 = ~(sub_718_2_n_95 | sub_718_2_n_74);
 assign sub_718_2_n_130 = ~(sub_718_2_n_9 & sub_718_2_n_77);
 assign sub_718_2_n_122 = ~(sub_718_2_n_93 | sub_718_2_n_49);
 assign sub_718_2_n_121 = ~(sub_718_2_n_97 | sub_718_2_n_80);
 assign sub_718_2_n_120 = ~(sub_718_2_n_65 | sub_718_2_n_89);
 assign sub_718_2_n_119 = ~(sub_718_2_n_76 | sub_718_2_n_94);
 assign sub_718_2_n_118 = ~(sub_718_2_n_90 | sub_718_2_n_78);
 assign sub_718_2_n_117 = ~(sub_718_2_n_79 | sub_718_2_n_69);
 assign sub_718_2_n_129 = ~(sub_718_2_n_85 | sub_718_2_n_51);
 assign sub_718_2_n_128 = ~(sub_718_2_n_5 | sub_718_2_n_74);
 assign sub_718_2_n_127 = ~(sub_718_2_n_99 | sub_718_2_n_94);
 assign sub_718_2_n_125 = ~(sub_718_2_n_6 | sub_718_2_n_80);
 assign sub_718_2_n_124 = ~(sub_718_2_n_83 | sub_718_2_n_50);
 assign sub_718_2_n_116 = ~(sub_718_2_n_82 | sub_718_2_n_87);
 assign in1_76_0_ = ~(sub_718_2_n_64 & ~(sub_718_2_n_57 & n_1542));
 assign sub_718_2_n_115 = ~(sub_718_2_n_88 | sub_718_2_n_80);
 assign sub_718_2_n_107 = ~(sub_718_2_n_98 | sub_718_2_n_89);
 assign sub_718_2_n_114 = ~(sub_718_2_n_1 | ~sub_718_2_n_101);
 assign sub_718_2_n_113 = ~(sub_718_2_n_10 | sub_718_2_n_94);
 assign sub_718_2_n_112 = ~(sub_718_2_n_81 | ~sub_718_2_n_103);
 assign sub_718_2_n_106 = ~(sub_718_2_n_102 | sub_718_2_n_69);
 assign sub_718_2_n_111 = ~(sub_718_2_n_84 | sub_718_2_n_49);
 assign sub_718_2_n_110 = ~(sub_718_2_n_100 | sub_718_2_n_74);
 assign sub_718_2_n_109 = ~(sub_718_2_n_86 | sub_718_2_n_78);
 assign sub_718_2_n_105 = ~(sub_718_2_n_92 & ~sub_718_2_n_75);
 assign sub_718_2_n_104 = ~(sub_718_2_n_95 & ~sub_718_2_n_5);
 assign sub_718_2_n_91 = ~sub_718_2_n_90;
 assign sub_718_2_n_103 = ~(in1_74_2_ & ~n_1579);
 assign sub_718_2_n_102 = (sub_718_2_n_58 & in1_74_18_);
 assign sub_718_2_n_101 = ~(in1_74_10_ & ~n_1555);
 assign sub_718_2_n_100 = (sub_718_2_n_60 & in1_74_12_);
 assign sub_718_2_n_99 = (sub_718_2_n_61 & in1_74_8_);
 assign sub_718_2_n_98 = (sub_718_2_n_55 & in1_74_16_);
 assign sub_718_2_n_97 = ~(in1_74_13_ & ~n_1577);
 assign sub_718_2_n_51 = ~(in1_74_22_ | sub_718_2_n_52);
 assign sub_718_2_n_96 = ~(in1_74_5_ | ~n_1567);
 assign sub_718_2_n_95 = ~(in1_74_11_ & ~n_1595);
 assign sub_718_2_n_94 = ~(in1_74_8_ | sub_718_2_n_61);
 assign sub_718_2_n_93 = ~(in1_74_5_ & ~n_1567);
 assign sub_718_2_n_92 = ~(in1_74_9_ & ~n_1551);
 assign sub_718_2_n_90 = ~(in1_74_3_ & ~n_1535);
 assign sub_718_2_n_89 = ~(in1_74_16_ | sub_718_2_n_55);
 assign sub_718_2_n_50 = ~(in1_74_20_ | sub_718_2_n_53);
 assign sub_718_2_n_49 = ~(in1_74_6_ | sub_718_2_n_56);
 assign sub_718_2_n_77 = ~sub_718_2_n_78;
 assign sub_718_2_n_73 = ~sub_718_2_n_72;
 assign sub_718_2_n_71 = ~sub_718_2_n_70;
 assign sub_718_2_n_68 = ~sub_718_2_n_67;
 assign sub_718_2_n_66 = ~sub_718_2_n_65;
 assign sub_718_2_n_88 = (sub_718_2_n_62 & in1_74_14_);
 assign sub_718_2_n_87 = ~(in1_74_0_ | sub_718_2_n_63);
 assign sub_718_2_n_86 = (sub_718_2_n_54 & in1_74_4_);
 assign sub_718_2_n_85 = (sub_718_2_n_52 & in1_74_22_);
 assign sub_718_2_n_84 = (sub_718_2_n_56 & in1_74_6_);
 assign sub_718_2_n_83 = (sub_718_2_n_53 & in1_74_20_);
 assign sub_718_2_n_82 = (sub_718_2_n_63 & in1_74_0_);
 assign sub_718_2_n_81 = ~(in1_74_2_ | sub_718_2_n_59);
 assign sub_718_2_n_80 = ~(in1_74_14_ | sub_718_2_n_62);
 assign sub_718_2_n_79 = ~(in1_74_17_ & ~n_1472);
 assign sub_718_2_n_78 = ~(in1_74_4_ | sub_718_2_n_54);
 assign sub_718_2_n_76 = ~(in1_74_7_ & ~n_1479);
 assign sub_718_2_n_75 = ~(in1_74_9_ | ~n_1551);
 assign sub_718_2_n_74 = ~(in1_74_12_ | sub_718_2_n_60);
 assign sub_718_2_n_72 = ~(in1_74_21_ & ~n_1591);
 assign sub_718_2_n_70 = ~(in1_74_19_ & ~n_1565);
 assign sub_718_2_n_69 = ~(in1_74_18_ | sub_718_2_n_58);
 assign sub_718_2_n_67 = ~(in1_74_1_ & ~n_1477);
 assign sub_718_2_n_65 = ~(in1_74_15_ & ~n_1549);
 assign sub_718_2_n_64 = ~(n_1543 & ~n_1542);
 assign sub_718_2_n_63 = ~n_1586;
 assign sub_718_2_n_62 = ~n_1495;
 assign sub_718_2_n_61 = ~n_1589;
 assign sub_718_2_n_60 = ~n_1581;
 assign sub_718_2_n_59 = ~n_1579;
 assign sub_718_2_n_58 = ~n_1558;
 assign sub_718_2_n_57 = ~n_1543;
 assign sub_718_2_n_56 = ~n_1527;
 assign sub_718_2_n_55 = ~n_1562;
 assign sub_718_2_n_54 = ~n_1569;
 assign sub_718_2_n_53 = ~n_1593;
 assign sub_718_2_n_52 = ~n_1403;
 assign in1_76_14_ = ~(sub_718_2_n_193 ^ sub_718_2_n_26);
 assign in1_76_10_ = (sub_718_2_n_178 ^ sub_718_2_n_105);
 assign sub_718_2_n_46 = ~(sub_718_2_n_174 | ~sub_718_2_n_163);
 assign in1_76_1_ = (sub_718_2_n_116 ^ sub_718_2_n_64);
 assign sub_718_2_n_44 = ~(sub_718_2_n_33 & ~sub_718_2_n_149);
 assign sub_718_2_n_43 = ~(sub_718_2_n_46 | ~sub_718_2_n_146);
 assign sub_718_2_n_42 = ~(sub_718_2_n_184 | ~sub_718_2_n_137);
 assign in1_76_23_ = ~(sub_718_2_n_202 ^ sub_718_2_n_129);
 assign in1_76_9_ = (sub_718_2_n_177 ^ sub_718_2_n_127);
 assign in1_76_6_ = ~(sub_718_2_n_170 ^ sub_718_2_n_23);
 assign in1_76_22_ = (sub_718_2_n_200 ^ sub_718_2_n_22);
 assign in1_76_21_ = ~(sub_718_2_n_199 ^ sub_718_2_n_124);
 assign in1_76_15_ = (sub_718_2_n_197 ^ sub_718_2_n_115);
 assign in1_76_4_ = ~(sub_718_2_n_166 ^ sub_718_2_n_16);
 assign in1_76_11_ = (sub_718_2_n_185 ^ sub_718_2_n_114);
 assign sub_718_2_n_33 = ~(sub_718_2_n_17 | ~sub_718_2_n_113);
 assign in1_76_3_ = ~(sub_718_2_n_167 ^ sub_718_2_n_112);
 assign in1_76_7_ = (sub_718_2_n_175 ^ sub_718_2_n_111);
 assign in1_76_13_ = (sub_718_2_n_186 ^ sub_718_2_n_110);
 assign in1_76_5_ = ~(sub_718_2_n_169 ^ sub_718_2_n_109);
 assign in1_76_20_ = (sub_718_2_n_192 ^ sub_718_2_n_24);
 assign in1_76_2_ = (sub_718_2_n_161 ^ sub_718_2_n_11);
 assign sub_718_2_n_26 = ~(sub_718_2_n_6 | ~sub_718_2_n_97);
 assign sub_718_2_n_25 = ~(sub_718_2_n_7 & ~sub_718_2_n_51);
 assign sub_718_2_n_24 = ~(sub_718_2_n_71 | ~sub_718_2_n_3);
 assign sub_718_2_n_23 = ~(sub_718_2_n_96 | ~sub_718_2_n_93);
 assign sub_718_2_n_22 = ~(sub_718_2_n_73 | ~sub_718_2_n_7);
 assign sub_718_2_n_21 = ~(sub_718_2_n_4 & ~sub_718_2_n_89);
 assign sub_718_2_n_20 = ~(sub_718_2_n_3 & ~sub_718_2_n_50);
 assign sub_718_2_n_19 = (sub_718_2_n_49 | sub_718_2_n_96);
 assign sub_718_2_n_18 = ~(sub_718_2_n_0 & ~sub_718_2_n_81);
 assign sub_718_2_n_17 = (sub_718_2_n_1 | sub_718_2_n_75);
 assign sub_718_2_n_16 = ~(sub_718_2_n_91 | ~sub_718_2_n_9);
 assign sub_718_2_n_15 = ~(sub_718_2_n_8 | ~sub_718_2_n_79);
 assign sub_718_2_n_14 = ~(sub_718_2_n_10 | ~sub_718_2_n_76);
 assign sub_718_2_n_13 = ~(sub_718_2_n_66 | ~sub_718_2_n_4);
 assign sub_718_2_n_12 = (sub_718_2_n_69 | sub_718_2_n_8);
 assign sub_718_2_n_11 = ~(sub_718_2_n_68 | ~sub_718_2_n_0);
 assign sub_718_2_n_10 = ~(in1_74_7_ | ~n_1479);
 assign sub_718_2_n_9 = ~(n_1535 & ~in1_74_3_);
 assign sub_718_2_n_8 = ~(in1_74_17_ | ~n_1472);
 assign sub_718_2_n_7 = ~(n_1591 & ~in1_74_21_);
 assign sub_718_2_n_6 = ~(in1_74_13_ | ~n_1577);
 assign sub_718_2_n_5 = ~(in1_74_11_ | ~n_1595);
 assign sub_718_2_n_4 = ~(n_1549 & ~in1_74_15_);
 assign sub_718_2_n_3 = ~(n_1565 & ~in1_74_19_);
 assign sub_718_2_n_2 = ~(sub_718_2_n_182 & ~in1_74_23_);
 assign sub_718_2_n_1 = ~(in1_74_10_ | ~n_1555);
 assign sub_718_2_n_0 = ~(n_1477 & ~in1_74_1_);
 assign sub_739_2_n_180 = ~(sub_739_2_n_67 & (sub_739_2_n_179 | sub_739_2_n_12));
 assign sub_739_2_n_179 = ~sub_739_2_n_178;
 assign sub_739_2_n_178 = ~(sub_739_2_n_121 & (sub_739_2_n_51 | sub_739_2_n_104));
 assign sub_739_2_n_177 = ~(sub_739_2_n_63 & (sub_739_2_n_51 | sub_739_2_n_82));
 assign sub_739_2_n_176 = ~(sub_739_2_n_83 & (sub_739_2_n_171 | sub_739_2_n_4));
 assign in1_79_20_ = ~(sub_739_2_n_51 ^ sub_739_2_n_16);
 assign in1_79_18_ = ~(sub_739_2_n_171 ^ sub_739_2_n_27);
 assign sub_739_2_n_173 = ~(sub_739_2_n_85 & (sub_739_2_n_166 | sub_739_2_n_73));
 assign in1_79_24_ = ~(sub_739_2_n_2 & sub_739_2_n_54);
 assign sub_739_2_n_171 = ~(sub_739_2_n_43 | sub_739_2_n_120);
 assign sub_739_2_n_170 = ~(sub_739_2_n_65 & (sub_739_2_n_53 | sub_739_2_n_13));
 assign in1_79_16_ = ~(sub_739_2_n_53 ^ sub_739_2_n_17);
 assign sub_739_2_n_168 = ~(sub_739_2_n_53 | sub_739_2_n_125);
 assign sub_739_2_n_167 = ~(sub_739_2_n_152 | ~(sub_739_2_n_161 | sub_739_2_n_50));
 assign sub_739_2_n_166 = ~sub_739_2_n_165;
 assign sub_739_2_n_165 = ~(sub_739_2_n_119 & (sub_739_2_n_160 | sub_739_2_n_29));
 assign sub_739_2_n_164 = ~(sub_739_2_n_81 & (sub_739_2_n_160 | sub_739_2_n_70));
 assign sub_739_2_n_163 = ~(sub_739_2_n_88 & (sub_739_2_n_159 | sub_739_2_n_11));
 assign in1_79_12_ = ~(sub_739_2_n_160 ^ sub_739_2_n_26);
 assign sub_739_2_n_161 = ~(sub_739_2_n_56 & (sub_739_2_n_128 & sub_739_2_n_126));
 assign sub_739_2_n_160 = ~(sub_739_2_n_139 | (sub_739_2_n_56 & sub_739_2_n_128));
 assign sub_739_2_n_159 = ~(sub_739_2_n_33 | sub_739_2_n_117);
 assign sub_739_2_n_158 = ~(sub_739_2_n_79 & (sub_739_2_n_156 | sub_739_2_n_69));
 assign sub_739_2_n_157 = ~(sub_739_2_n_80 & (sub_739_2_n_49 | sub_739_2_n_3));
 assign sub_739_2_n_156 = ~sub_739_2_n_56;
 assign sub_739_2_n_56 = ~(sub_739_2_n_138 & (sub_739_2_n_148 | (sub_739_2_n_19 | sub_739_2_n_22)));
 assign sub_739_2_n_155 = ~(sub_739_2_n_87 | (sub_739_2_n_147 & sub_739_2_n_1));
 assign in1_79_4_ = ~(sub_739_2_n_147 ^ sub_739_2_n_105);
 assign in1_79_3_ = (sub_739_2_n_150 ^ sub_739_2_n_95);
 assign sub_739_2_n_152 = ~(sub_739_2_n_151 & sub_739_2_n_143);
 assign sub_739_2_n_151 = ~(sub_739_2_n_144 & ~sub_739_2_n_50);
 assign sub_739_2_n_150 = ~(sub_739_2_n_84 & (sub_739_2_n_142 | sub_739_2_n_66));
 assign in1_79_2_ = ~(sub_739_2_n_146 & ~sub_739_2_n_145);
 assign sub_739_2_n_147 = ~sub_739_2_n_148;
 assign sub_739_2_n_148 = ~(sub_739_2_n_116 | (sub_739_2_n_135 & sub_739_2_n_97));
 assign sub_739_2_n_146 = ~(sub_739_2_n_135 & sub_739_2_n_113);
 assign sub_739_2_n_145 = ~(sub_739_2_n_135 | sub_739_2_n_113);
 assign sub_739_2_n_144 = ~(sub_739_2_n_137 & ~(sub_739_2_n_139 & sub_739_2_n_126));
 assign sub_739_2_n_143 = ~(sub_739_2_n_141 | sub_739_2_n_136);
 assign sub_739_2_n_142 = ~sub_739_2_n_135;
 assign sub_739_2_n_141 = ~(sub_739_2_n_140 | sub_739_2_n_127);
 assign sub_739_2_n_140 = ~(sub_739_2_n_122 | (sub_739_2_n_120 & sub_739_2_n_108));
 assign sub_739_2_n_139 = ~(sub_739_2_n_133 & sub_739_2_n_115);
 assign sub_739_2_n_138 = ~(sub_739_2_n_132 | sub_739_2_n_123);
 assign sub_739_2_n_137 = ~(sub_739_2_n_124 | ~(sub_739_2_n_119 | sub_739_2_n_24));
 assign sub_739_2_n_136 = ~(sub_739_2_n_130 & sub_739_2_n_114);
 assign sub_739_2_n_135 = ~(sub_739_2_n_131 & sub_739_2_n_90);
 assign in1_79_1_ = ~((sub_739_2_n_129 & ~sub_739_2_n_32) | (sub_739_2_n_62 & sub_739_2_n_32));
 assign sub_739_2_n_133 = ~(sub_739_2_n_117 & sub_739_2_n_103);
 assign sub_739_2_n_132 = ~(sub_739_2_n_118 | sub_739_2_n_22);
 assign sub_739_2_n_131 = ~(sub_739_2_n_14 & ~sub_739_2_n_129);
 assign sub_739_2_n_130 = ~(sub_739_2_n_111 & ~sub_739_2_n_121);
 assign sub_739_2_n_129 = ~sub_739_2_n_62;
 assign sub_739_2_n_124 = ~(sub_739_2_n_76 & (sub_739_2_n_85 | sub_739_2_n_9));
 assign sub_739_2_n_123 = ~(sub_739_2_n_89 & (sub_739_2_n_80 | sub_739_2_n_10));
 assign sub_739_2_n_128 = (sub_739_2_n_98 & sub_739_2_n_103);
 assign sub_739_2_n_122 = ~(sub_739_2_n_77 & (sub_739_2_n_83 | sub_739_2_n_0));
 assign sub_739_2_n_127 = ~(sub_739_2_n_111 & ~sub_739_2_n_104);
 assign sub_739_2_n_126 = ~(sub_739_2_n_29 | sub_739_2_n_24);
 assign sub_739_2_n_125 = ~(sub_739_2_n_107 & sub_739_2_n_108);
 assign sub_739_2_n_116 = ~(sub_739_2_n_91 & (sub_739_2_n_84 | sub_739_2_n_6));
 assign sub_739_2_n_115 = ~(sub_739_2_n_93 | ~(sub_739_2_n_88 | sub_739_2_n_64));
 assign sub_739_2_n_114 = ~(sub_739_2_n_78 | ~(sub_739_2_n_67 | sub_739_2_n_71));
 assign sub_739_2_n_121 = ~(sub_739_2_n_15 | ~(sub_739_2_n_63 | sub_739_2_n_72));
 assign sub_739_2_n_120 = ~(sub_739_2_n_75 & (sub_739_2_n_65 | sub_739_2_n_5));
 assign sub_739_2_n_119 = ~(sub_739_2_n_94 | ~(sub_739_2_n_81 | sub_739_2_n_55));
 assign sub_739_2_n_118 = ~(sub_739_2_n_106 | sub_739_2_n_92);
 assign sub_739_2_n_117 = ~(sub_739_2_n_74 & (sub_739_2_n_79 | sub_739_2_n_8));
 assign sub_739_2_n_106 = ~(sub_739_2_n_86 | sub_739_2_n_68);
 assign sub_739_2_n_113 = ~(sub_739_2_n_84 & ~sub_739_2_n_66);
 assign sub_739_2_n_112 = ~(sub_739_2_n_78 | sub_739_2_n_71);
 assign sub_739_2_n_105 = ~(sub_739_2_n_86 & sub_739_2_n_1);
 assign sub_739_2_n_111 = ~(sub_739_2_n_12 | sub_739_2_n_71);
 assign sub_739_2_n_110 = ~(sub_739_2_n_92 | sub_739_2_n_68);
 assign sub_739_2_n_109 = ~(sub_739_2_n_15 | sub_739_2_n_72);
 assign sub_739_2_n_108 = ~(sub_739_2_n_4 | sub_739_2_n_0);
 assign sub_739_2_n_107 = ~(sub_739_2_n_13 | sub_739_2_n_5);
 assign sub_739_2_n_97 = ~(sub_739_2_n_66 | sub_739_2_n_6);
 assign in1_79_0_ = ~(sub_739_2_n_62 & ~(sub_739_2_n_60 & n_1585));
 assign sub_739_2_n_104 = (sub_739_2_n_82 | sub_739_2_n_72);
 assign sub_739_2_n_95 = ~(sub_739_2_n_6 | ~sub_739_2_n_91);
 assign sub_739_2_n_103 = ~(sub_739_2_n_11 | sub_739_2_n_64);
 assign sub_739_2_n_102 = ~(sub_739_2_n_0 | ~sub_739_2_n_77);
 assign sub_739_2_n_101 = ~(sub_739_2_n_94 | sub_739_2_n_55);
 assign sub_739_2_n_100 = ~(sub_739_2_n_93 | sub_739_2_n_64);
 assign sub_739_2_n_99 = ~(sub_739_2_n_9 | ~sub_739_2_n_76);
 assign sub_739_2_n_98 = ~(sub_739_2_n_69 | sub_739_2_n_8);
 assign sub_739_2_n_87 = ~sub_739_2_n_86;
 assign sub_739_2_n_94 = (sub_739_2_n_57 & in1_77_12_);
 assign sub_739_2_n_93 = (sub_739_2_n_58 & in1_77_10_);
 assign sub_739_2_n_92 = (sub_739_2_n_61 & in1_77_4_);
 assign sub_739_2_n_91 = ~(in1_77_2_ & ~n_1579);
 assign sub_739_2_n_90 = ~(in1_77_0_ & ~n_1586);
 assign sub_739_2_n_89 = ~(in1_77_6_ & ~n_1527);
 assign sub_739_2_n_88 = ~(in1_77_9_ & ~n_1551);
 assign sub_739_2_n_55 = ~(in1_77_12_ | sub_739_2_n_57);
 assign sub_739_2_n_86 = ~(in1_77_3_ & ~n_1535);
 assign sub_739_2_n_85 = ~(in1_77_13_ & ~n_1577);
 assign sub_739_2_n_84 = ~(in1_77_1_ & ~n_1477);
 assign sub_739_2_n_83 = ~(in1_77_17_ & ~n_1472);
 assign sub_739_2_n_82 = ~(in1_77_19_ | ~n_1565);
 assign sub_739_2_n_81 = ~(in1_77_11_ & ~n_1595);
 assign sub_739_2_n_80 = ~(in1_77_5_ & ~n_1567);
 assign sub_739_2_n_79 = ~(in1_77_7_ & ~n_1479);
 assign sub_739_2_n_70 = ~sub_739_2_n_7;
 assign sub_739_2_n_78 = (sub_739_2_n_59 & in1_77_22_);
 assign sub_739_2_n_77 = ~(in1_77_18_ & ~n_1558);
 assign sub_739_2_n_76 = ~(in1_77_14_ & ~n_1495);
 assign sub_739_2_n_75 = ~(in1_77_16_ & ~n_1562);
 assign sub_739_2_n_74 = ~(in1_77_8_ & ~n_1589);
 assign sub_739_2_n_73 = ~(in1_77_13_ | ~n_1577);
 assign sub_739_2_n_72 = ~(in1_77_20_ | ~n_1593);
 assign sub_739_2_n_71 = ~(in1_77_22_ | sub_739_2_n_59);
 assign sub_739_2_n_69 = ~(in1_77_7_ | ~n_1479);
 assign sub_739_2_n_68 = ~(in1_77_4_ | sub_739_2_n_61);
 assign sub_739_2_n_67 = ~(in1_77_21_ & ~n_1591);
 assign sub_739_2_n_66 = ~(in1_77_1_ | ~n_1477);
 assign sub_739_2_n_65 = ~(in1_77_15_ & ~n_1549);
 assign sub_739_2_n_64 = ~(in1_77_10_ | sub_739_2_n_58);
 assign sub_739_2_n_63 = ~(in1_77_19_ & ~n_1565);
 assign sub_739_2_n_62 = ~(n_1543 & ~n_1585);
 assign sub_739_2_n_61 = ~n_1569;
 assign sub_739_2_n_60 = ~n_1543;
 assign sub_739_2_n_59 = ~n_1403;
 assign sub_739_2_n_58 = ~n_1555;
 assign sub_739_2_n_57 = ~n_1581;
 assign sub_739_2_n_54 = ~(in1_77_23_ & ~sub_739_2_n_167);
 assign sub_739_2_n_53 = ~(sub_739_2_n_144 | ~sub_739_2_n_161);
 assign in1_79_10_ = ~(sub_739_2_n_159 ^ sub_739_2_n_30);
 assign sub_739_2_n_51 = ~(sub_739_2_n_168 | ~sub_739_2_n_140);
 assign sub_739_2_n_50 = (sub_739_2_n_127 | sub_739_2_n_125);
 assign sub_739_2_n_49 = (sub_739_2_n_118 & (sub_739_2_n_148 | sub_739_2_n_19));
 assign in1_79_23_ = (sub_739_2_n_180 ^ sub_739_2_n_112);
 assign in1_79_9_ = (sub_739_2_n_158 ^ sub_739_2_n_20);
 assign in1_79_5_ = ~(sub_739_2_n_155 ^ sub_739_2_n_110);
 assign in1_79_22_ = (sub_739_2_n_178 ^ sub_739_2_n_18);
 assign in1_79_21_ = (sub_739_2_n_177 ^ sub_739_2_n_109);
 assign sub_739_2_n_43 = ~(sub_739_2_n_53 | ~sub_739_2_n_107);
 assign in1_79_17_ = (sub_739_2_n_170 ^ sub_739_2_n_21);
 assign in1_79_6_ = ~(sub_739_2_n_49 ^ sub_739_2_n_25);
 assign in1_79_7_ = (sub_739_2_n_157 ^ sub_739_2_n_31);
 assign in1_79_19_ = (sub_739_2_n_176 ^ sub_739_2_n_102);
 assign in1_79_14_ = (sub_739_2_n_165 ^ sub_739_2_n_28);
 assign in1_79_13_ = (sub_739_2_n_164 ^ sub_739_2_n_101);
 assign in1_79_8_ = (sub_739_2_n_56 ^ sub_739_2_n_23);
 assign in1_79_11_ = (sub_739_2_n_163 ^ sub_739_2_n_100);
 assign in1_79_15_ = (sub_739_2_n_173 ^ sub_739_2_n_99);
 assign sub_739_2_n_33 = ~(sub_739_2_n_156 | ~sub_739_2_n_98);
 assign sub_739_2_n_32 = (sub_739_2_n_90 & sub_739_2_n_14);
 assign sub_739_2_n_31 = ~(sub_739_2_n_10 | ~sub_739_2_n_89);
 assign sub_739_2_n_30 = ~(sub_739_2_n_11 | ~sub_739_2_n_88);
 assign sub_739_2_n_29 = ~(sub_739_2_n_7 & ~sub_739_2_n_55);
 assign sub_739_2_n_28 = ~(sub_739_2_n_73 | ~sub_739_2_n_85);
 assign sub_739_2_n_27 = ~(sub_739_2_n_4 | ~sub_739_2_n_83);
 assign sub_739_2_n_26 = ~(sub_739_2_n_70 | ~sub_739_2_n_81);
 assign sub_739_2_n_25 = ~(sub_739_2_n_3 | ~sub_739_2_n_80);
 assign sub_739_2_n_24 = (sub_739_2_n_9 | sub_739_2_n_73);
 assign sub_739_2_n_23 = ~(sub_739_2_n_69 | ~sub_739_2_n_79);
 assign sub_739_2_n_22 = (sub_739_2_n_10 | sub_739_2_n_3);
 assign sub_739_2_n_21 = ~(sub_739_2_n_5 | ~sub_739_2_n_75);
 assign sub_739_2_n_20 = ~(sub_739_2_n_8 | ~sub_739_2_n_74);
 assign sub_739_2_n_19 = ~(sub_739_2_n_1 & ~sub_739_2_n_68);
 assign sub_739_2_n_18 = ~(sub_739_2_n_12 | ~sub_739_2_n_67);
 assign sub_739_2_n_17 = ~(sub_739_2_n_13 | ~sub_739_2_n_65);
 assign sub_739_2_n_16 = ~(sub_739_2_n_82 | ~sub_739_2_n_63);
 assign sub_739_2_n_15 = ~(n_1593 | ~in1_77_20_);
 assign sub_739_2_n_14 = ~(n_1586 & ~in1_77_0_);
 assign sub_739_2_n_13 = ~(in1_77_15_ | ~n_1549);
 assign sub_739_2_n_12 = ~(in1_77_21_ | ~n_1591);
 assign sub_739_2_n_11 = ~(in1_77_9_ | ~n_1551);
 assign sub_739_2_n_10 = ~(in1_77_6_ | ~n_1527);
 assign sub_739_2_n_9 = ~(in1_77_14_ | ~n_1495);
 assign sub_739_2_n_8 = ~(in1_77_8_ | ~n_1589);
 assign sub_739_2_n_7 = ~(n_1595 & ~in1_77_11_);
 assign sub_739_2_n_6 = ~(in1_77_2_ | ~n_1579);
 assign sub_739_2_n_5 = ~(in1_77_16_ | ~n_1562);
 assign sub_739_2_n_4 = ~(in1_77_17_ | ~n_1472);
 assign sub_739_2_n_3 = ~(in1_77_5_ | ~n_1567);
 assign sub_739_2_n_2 = ~(sub_739_2_n_167 & ~in1_77_23_);
 assign sub_739_2_n_1 = ~(n_1535 & ~in1_77_3_);
 assign sub_739_2_n_0 = ~(in1_77_18_ | ~n_1558);
 assign sub_760_2_n_174 = ~(sub_760_2_n_63 & (sub_760_2_n_172 | sub_760_2_n_79));
 assign in1_82_21_ = (sub_760_2_n_171 ^ sub_760_2_n_21);
 assign sub_760_2_n_172 = ~(sub_760_2_n_115 | (sub_760_2_n_163 & sub_760_2_n_97));
 assign sub_760_2_n_171 = ~(sub_760_2_n_62 & (sub_760_2_n_164 | sub_760_2_n_4));
 assign sub_760_2_n_170 = ~(sub_760_2_n_67 & (sub_760_2_n_165 | sub_760_2_n_13));
 assign sub_760_2_n_169 = ~(sub_760_2_n_86 & (sub_760_2_n_166 | sub_760_2_n_10));
 assign in1_82_18_ = ~(sub_760_2_n_165 ^ sub_760_2_n_19);
 assign in1_82_24_ = ~(sub_760_2_n_162 & sub_760_2_n_161);
 assign sub_760_2_n_164 = ~sub_760_2_n_163;
 assign sub_760_2_n_162 = ~(sub_760_2_n_156 & sub_760_2_n_56);
 assign sub_760_2_n_161 = ~(sub_760_2_n_155 & in1_80_23_);
 assign sub_760_2_n_160 = ~(sub_760_2_n_59 & (sub_760_2_n_153 | sub_760_2_n_64));
 assign sub_760_2_n_166 = ~(sub_760_2_n_116 | (sub_760_2_n_152 & sub_760_2_n_102));
 assign sub_760_2_n_165 = ~(sub_760_2_n_34 | sub_760_2_n_114);
 assign sub_760_2_n_163 = ~(sub_760_2_n_129 & (sub_760_2_n_153 | sub_760_2_n_121));
 assign in1_82_16_ = ~(sub_760_2_n_153 ^ sub_760_2_n_14);
 assign sub_760_2_n_158 = ~(sub_760_2_n_85 & ~(sub_760_2_n_152 & sub_760_2_n_80));
 assign sub_760_2_n_157 = ~(sub_760_2_n_81 & (sub_760_2_n_151 | sub_760_2_n_65));
 assign sub_760_2_n_156 = ~sub_760_2_n_155;
 assign sub_760_2_n_155 = ~(sub_760_2_n_140 & sub_760_2_n_154);
 assign sub_760_2_n_154 = ~(sub_760_2_n_146 & sub_760_2_n_126);
 assign sub_760_2_n_153 = ~(sub_760_2_n_146 | sub_760_2_n_134);
 assign sub_760_2_n_152 = ~(sub_760_2_n_148 & sub_760_2_n_132);
 assign sub_760_2_n_151 = ~sub_760_2_n_150;
 assign sub_760_2_n_150 = ~(sub_760_2_n_113 & (sub_760_2_n_145 | sub_760_2_n_98));
 assign sub_760_2_n_149 = ~(sub_760_2_n_66 & (sub_760_2_n_145 | sub_760_2_n_83));
 assign sub_760_2_n_148 = ~(sub_760_2_n_144 & sub_760_2_n_123);
 assign sub_760_2_n_147 = ~(sub_760_2_n_82 & (sub_760_2_n_143 | sub_760_2_n_2));
 assign sub_760_2_n_146 = ~(sub_760_2_n_145 | sub_760_2_n_52);
 assign sub_760_2_n_144 = ~sub_760_2_n_145;
 assign sub_760_2_n_145 = ~(sub_760_2_n_48 | sub_760_2_n_131);
 assign sub_760_2_n_143 = ~(sub_760_2_n_117 | ~(sub_760_2_n_136 | sub_760_2_n_109));
 assign sub_760_2_n_142 = ~(sub_760_2_n_78 & (sub_760_2_n_136 | sub_760_2_n_68));
 assign in1_82_3_ = (sub_760_2_n_138 ^ sub_760_2_n_93);
 assign sub_760_2_n_140 = ~(sub_760_2_n_139 | sub_760_2_n_133);
 assign sub_760_2_n_139 = (sub_760_2_n_134 & sub_760_2_n_126);
 assign sub_760_2_n_138 = ~(sub_760_2_n_61 & (sub_760_2_n_127 | sub_760_2_n_60));
 assign in1_82_2_ = ~(sub_760_2_n_127 ^ sub_760_2_n_15);
 assign sub_760_2_n_136 = ~(sub_760_2_n_135 | sub_760_2_n_111);
 assign sub_760_2_n_135 = ~(sub_760_2_n_127 | sub_760_2_n_20);
 assign sub_760_2_n_134 = ~(sub_760_2_n_130 & (sub_760_2_n_132 | sub_760_2_n_124));
 assign sub_760_2_n_133 = ~(sub_760_2_n_51 & sub_760_2_n_128);
 assign sub_760_2_n_132 = ~(sub_760_2_n_112 | ~(sub_760_2_n_113 | sub_760_2_n_99));
 assign sub_760_2_n_131 = ~(sub_760_2_n_119 & ~(sub_760_2_n_117 & sub_760_2_n_107));
 assign sub_760_2_n_130 = ~(sub_760_2_n_120 | (sub_760_2_n_116 & sub_760_2_n_105));
 assign sub_760_2_n_129 = ~(sub_760_2_n_118 | (sub_760_2_n_114 & sub_760_2_n_103));
 assign sub_760_2_n_128 = ~(sub_760_2_n_45 | sub_760_2_n_110);
 assign sub_760_2_n_127 = ~(sub_760_2_n_125 | sub_760_2_n_7);
 assign sub_760_2_n_126 = ~(sub_760_2_n_121 | sub_760_2_n_122);
 assign sub_760_2_n_125 = ~(sub_760_2_n_75 | ~sub_760_2_n_58);
 assign sub_760_2_n_120 = ~(sub_760_2_n_76 & (sub_760_2_n_86 | sub_760_2_n_12));
 assign sub_760_2_n_119 = ~(sub_760_2_n_72 | ~(sub_760_2_n_82 | sub_760_2_n_77));
 assign sub_760_2_n_118 = ~(sub_760_2_n_91 & (sub_760_2_n_67 | sub_760_2_n_8));
 assign sub_760_2_n_124 = ~(sub_760_2_n_102 & sub_760_2_n_105);
 assign sub_760_2_n_123 = ~(sub_760_2_n_98 | sub_760_2_n_99);
 assign sub_760_2_n_122 = ~(sub_760_2_n_97 & sub_760_2_n_104);
 assign sub_760_2_n_121 = ~(sub_760_2_n_95 & sub_760_2_n_103);
 assign sub_760_2_n_112 = ~(sub_760_2_n_90 & (sub_760_2_n_81 | sub_760_2_n_1));
 assign sub_760_2_n_111 = ~(sub_760_2_n_92 & (sub_760_2_n_61 | sub_760_2_n_70));
 assign sub_760_2_n_110 = ~(sub_760_2_n_73 & (sub_760_2_n_63 | sub_760_2_n_0));
 assign sub_760_2_n_117 = ~(sub_760_2_n_74 & (sub_760_2_n_78 | sub_760_2_n_5));
 assign sub_760_2_n_116 = ~(sub_760_2_n_89 & (sub_760_2_n_85 | sub_760_2_n_11));
 assign sub_760_2_n_115 = ~(sub_760_2_n_71 & (sub_760_2_n_62 | sub_760_2_n_3));
 assign sub_760_2_n_114 = ~(sub_760_2_n_87 & (sub_760_2_n_59 | sub_760_2_n_6));
 assign sub_760_2_n_113 = ~(sub_760_2_n_88 | ~(sub_760_2_n_66 | sub_760_2_n_84));
 assign sub_760_2_n_109 = (sub_760_2_n_68 | sub_760_2_n_5);
 assign sub_760_2_n_101 = ~(sub_760_2_n_7 | sub_760_2_n_75);
 assign sub_760_2_n_108 = ~(sub_760_2_n_0 | ~sub_760_2_n_73);
 assign sub_760_2_n_107 = ~(sub_760_2_n_2 | sub_760_2_n_77);
 assign sub_760_2_n_106 = ~(sub_760_2_n_88 | sub_760_2_n_84);
 assign sub_760_2_n_105 = ~(sub_760_2_n_10 | sub_760_2_n_12);
 assign sub_760_2_n_104 = ~(sub_760_2_n_79 | sub_760_2_n_0);
 assign sub_760_2_n_103 = ~(sub_760_2_n_13 | sub_760_2_n_8);
 assign sub_760_2_n_102 = ~(sub_760_2_n_9 | sub_760_2_n_11);
 assign in1_82_0_ = ~(sub_760_2_n_58 & ~(sub_760_2_n_57 & n_1588));
 assign sub_760_2_n_100 = ~(sub_760_2_n_1 | ~sub_760_2_n_90);
 assign sub_760_2_n_99 = ~(sub_760_2_n_69 & ~sub_760_2_n_65);
 assign sub_760_2_n_98 = (sub_760_2_n_83 | sub_760_2_n_84);
 assign sub_760_2_n_93 = ~(sub_760_2_n_70 | ~sub_760_2_n_92);
 assign sub_760_2_n_97 = ~(sub_760_2_n_4 | sub_760_2_n_3);
 assign sub_760_2_n_96 = ~(sub_760_2_n_72 | sub_760_2_n_77);
 assign sub_760_2_n_95 = ~(sub_760_2_n_64 | sub_760_2_n_6);
 assign sub_760_2_n_80 = ~sub_760_2_n_9;
 assign sub_760_2_n_92 = ~(in1_80_2_ & ~n_1579);
 assign sub_760_2_n_91 = ~(in1_80_18_ & ~n_1558);
 assign sub_760_2_n_90 = ~(in1_80_10_ & ~n_1555);
 assign sub_760_2_n_89 = ~(in1_80_12_ & ~n_1581);
 assign sub_760_2_n_88 = ~(n_1589 | ~in1_80_8_);
 assign sub_760_2_n_87 = ~(in1_80_16_ & ~n_1562);
 assign sub_760_2_n_86 = ~(in1_80_13_ & ~n_1577);
 assign sub_760_2_n_85 = ~(in1_80_11_ & ~n_1595);
 assign sub_760_2_n_84 = ~(in1_80_8_ | ~n_1589);
 assign sub_760_2_n_83 = ~(in1_80_7_ | ~n_1479);
 assign sub_760_2_n_82 = ~(in1_80_5_ & ~n_1567);
 assign sub_760_2_n_81 = ~(in1_80_9_ & ~n_1551);
 assign sub_760_2_n_79 = ~(in1_80_21_ | sub_760_2_n_55);
 assign sub_760_2_n_78 = ~(in1_80_3_ & ~n_1535);
 assign sub_760_2_n_77 = ~(in1_80_6_ | ~n_1527);
 assign sub_760_2_n_69 = ~sub_760_2_n_1;
 assign sub_760_2_n_76 = ~(in1_80_14_ & ~n_1495);
 assign sub_760_2_n_75 = ~(in1_80_0_ | ~n_1586);
 assign sub_760_2_n_74 = ~(in1_80_4_ & ~n_1569);
 assign sub_760_2_n_73 = ~(in1_80_22_ & ~n_1403);
 assign sub_760_2_n_72 = ~(n_1527 | ~in1_80_6_);
 assign sub_760_2_n_71 = ~(in1_80_20_ & ~n_1593);
 assign sub_760_2_n_70 = ~(in1_80_2_ | ~n_1579);
 assign sub_760_2_n_68 = ~(in1_80_3_ | ~n_1535);
 assign sub_760_2_n_67 = ~(in1_80_17_ & ~n_1472);
 assign sub_760_2_n_66 = ~(in1_80_7_ & ~n_1479);
 assign sub_760_2_n_65 = ~(in1_80_9_ | ~n_1551);
 assign sub_760_2_n_64 = ~(in1_80_15_ | ~n_1549);
 assign sub_760_2_n_63 = ~(sub_760_2_n_55 & in1_80_21_);
 assign sub_760_2_n_62 = ~(in1_80_19_ & ~n_1565);
 assign sub_760_2_n_61 = ~(in1_80_1_ & ~n_1477);
 assign sub_760_2_n_60 = ~(in1_80_1_ | ~n_1477);
 assign sub_760_2_n_59 = ~(in1_80_15_ & ~n_1549);
 assign sub_760_2_n_58 = ~(n_1543 & ~n_1588);
 assign sub_760_2_n_57 = ~n_1543;
 assign sub_760_2_n_56 = ~in1_80_23_;
 assign sub_760_2_n_55 = ~n_1591;
 assign in1_82_14_ = ~(sub_760_2_n_166 ^ sub_760_2_n_28);
 assign in1_82_1_ = (sub_760_2_n_101 ^ sub_760_2_n_58);
 assign sub_760_2_n_52 = ~(sub_760_2_n_123 & ~sub_760_2_n_124);
 assign sub_760_2_n_51 = (sub_760_2_n_122 | sub_760_2_n_129);
 assign in1_82_8_ = (sub_760_2_n_144 ^ sub_760_2_n_18);
 assign in1_82_23_ = (sub_760_2_n_174 ^ sub_760_2_n_108);
 assign sub_760_2_n_48 = ~(sub_760_2_n_136 | (sub_760_2_n_109 | ~sub_760_2_n_107));
 assign in1_82_9_ = (sub_760_2_n_149 ^ sub_760_2_n_106);
 assign in1_82_6_ = ~(sub_760_2_n_143 ^ sub_760_2_n_26);
 assign sub_760_2_n_45 = (sub_760_2_n_104 & sub_760_2_n_115);
 assign in1_82_22_ = ~(sub_760_2_n_172 ^ sub_760_2_n_17);
 assign in1_82_20_ = (sub_760_2_n_163 ^ sub_760_2_n_16);
 assign in1_82_19_ = (sub_760_2_n_170 ^ sub_760_2_n_31);
 assign in1_82_4_ = ~(sub_760_2_n_136 ^ sub_760_2_n_24);
 assign in1_82_17_ = (sub_760_2_n_160 ^ sub_760_2_n_29);
 assign in1_82_11_ = (sub_760_2_n_157 ^ sub_760_2_n_100);
 assign in1_82_15_ = (sub_760_2_n_169 ^ sub_760_2_n_23);
 assign in1_82_7_ = (sub_760_2_n_147 ^ sub_760_2_n_96);
 assign in1_82_13_ = (sub_760_2_n_158 ^ sub_760_2_n_30);
 assign in1_82_5_ = (sub_760_2_n_142 ^ sub_760_2_n_22);
 assign sub_760_2_n_34 = ~(sub_760_2_n_153 | ~sub_760_2_n_95);
 assign in1_82_10_ = (sub_760_2_n_150 ^ sub_760_2_n_25);
 assign in1_82_12_ = (sub_760_2_n_152 ^ sub_760_2_n_27);
 assign sub_760_2_n_31 = ~(sub_760_2_n_8 | ~sub_760_2_n_91);
 assign sub_760_2_n_30 = ~(sub_760_2_n_11 | ~sub_760_2_n_89);
 assign sub_760_2_n_29 = ~(sub_760_2_n_6 | ~sub_760_2_n_87);
 assign sub_760_2_n_28 = ~(sub_760_2_n_10 | ~sub_760_2_n_86);
 assign sub_760_2_n_27 = ~(sub_760_2_n_9 | ~sub_760_2_n_85);
 assign sub_760_2_n_26 = ~(sub_760_2_n_2 | ~sub_760_2_n_82);
 assign sub_760_2_n_25 = ~(sub_760_2_n_65 | ~sub_760_2_n_81);
 assign sub_760_2_n_24 = ~(sub_760_2_n_68 | ~sub_760_2_n_78);
 assign sub_760_2_n_23 = ~(sub_760_2_n_12 | ~sub_760_2_n_76);
 assign sub_760_2_n_22 = ~(sub_760_2_n_5 | ~sub_760_2_n_74);
 assign sub_760_2_n_21 = ~(sub_760_2_n_3 | ~sub_760_2_n_71);
 assign sub_760_2_n_20 = (sub_760_2_n_70 | sub_760_2_n_60);
 assign sub_760_2_n_19 = ~(sub_760_2_n_13 | ~sub_760_2_n_67);
 assign sub_760_2_n_18 = ~(sub_760_2_n_83 | ~sub_760_2_n_66);
 assign sub_760_2_n_17 = ~(sub_760_2_n_79 | ~sub_760_2_n_63);
 assign sub_760_2_n_16 = ~(sub_760_2_n_4 | ~sub_760_2_n_62);
 assign sub_760_2_n_15 = ~(sub_760_2_n_60 | ~sub_760_2_n_61);
 assign sub_760_2_n_14 = ~(sub_760_2_n_64 | ~sub_760_2_n_59);
 assign sub_760_2_n_13 = ~(in1_80_17_ | ~n_1472);
 assign sub_760_2_n_12 = ~(in1_80_14_ | ~n_1495);
 assign sub_760_2_n_11 = ~(in1_80_12_ | ~n_1581);
 assign sub_760_2_n_10 = ~(in1_80_13_ | ~n_1577);
 assign sub_760_2_n_9 = ~(in1_80_11_ | ~n_1595);
 assign sub_760_2_n_8 = ~(in1_80_18_ | ~n_1558);
 assign sub_760_2_n_7 = ~(n_1586 | ~in1_80_0_);
 assign sub_760_2_n_6 = ~(in1_80_16_ | ~n_1562);
 assign sub_760_2_n_5 = ~(in1_80_4_ | ~n_1569);
 assign sub_760_2_n_4 = ~(in1_80_19_ | ~n_1565);
 assign sub_760_2_n_3 = ~(in1_80_20_ | ~n_1593);
 assign sub_760_2_n_2 = ~(in1_80_5_ | ~n_1567);
 assign sub_760_2_n_1 = ~(in1_80_10_ | ~n_1555);
 assign sub_760_2_n_0 = ~(in1_80_22_ | ~n_1403);
 assign sub_781_2_n_178 = ~(sub_781_2_n_46 | (sub_781_2_n_177 & sub_781_2_n_48));
 assign sub_781_2_n_177 = ~(sub_781_2_n_119 & (sub_781_2_n_169 | sub_781_2_n_96));
 assign sub_781_2_n_176 = ~(sub_781_2_n_67 & (sub_781_2_n_169 | sub_781_2_n_75));
 assign sub_781_2_n_175 = ~(sub_781_2_n_40 | (sub_781_2_n_168 & sub_781_2_n_57));
 assign sub_781_2_n_174 = ~(sub_781_2_n_51 & (sub_781_2_n_166 | sub_781_2_n_66));
 assign in1_85_14_ = (sub_781_2_n_166 ^ sub_781_2_n_87);
 assign in1_85_13_ = (sub_781_2_n_165 ^ sub_781_2_n_7);
 assign in1_85_11_ = (sub_781_2_n_164 ^ sub_781_2_n_86);
 assign in1_85_24_ = ((sub_781_2_n_36 & ~sub_781_2_n_161) | (in1_83_23_ & sub_781_2_n_161));
 assign sub_781_2_n_169 = ~(sub_781_2_n_162 | sub_781_2_n_137);
 assign sub_781_2_n_168 = ~(sub_781_2_n_120 & (sub_781_2_n_159 | sub_781_2_n_111));
 assign sub_781_2_n_167 = ~(sub_781_2_n_78 & (sub_781_2_n_159 | sub_781_2_n_52));
 assign sub_781_2_n_166 = ~(sub_781_2_n_125 | (sub_781_2_n_158 & sub_781_2_n_101));
 assign sub_781_2_n_165 = ~(sub_781_2_n_77 | (sub_781_2_n_158 & sub_781_2_n_55));
 assign sub_781_2_n_164 = ~(sub_781_2_n_72 | (sub_781_2_n_157 & sub_781_2_n_4));
 assign in1_85_16_ = ~(sub_781_2_n_159 ^ sub_781_2_n_14);
 assign sub_781_2_n_162 = ~(sub_781_2_n_159 | sub_781_2_n_128);
 assign sub_781_2_n_161 = ~(sub_781_2_n_147 & sub_781_2_n_160);
 assign sub_781_2_n_160 = ~(sub_781_2_n_154 & sub_781_2_n_129);
 assign sub_781_2_n_159 = ~(sub_781_2_n_154 | sub_781_2_n_143);
 assign sub_781_2_n_158 = ~(sub_781_2_n_135 & (sub_781_2_n_151 | sub_781_2_n_21));
 assign sub_781_2_n_157 = ~(sub_781_2_n_121 & (sub_781_2_n_151 | sub_781_2_n_107));
 assign sub_781_2_n_156 = ~(sub_781_2_n_39 & (sub_781_2_n_151 | sub_781_2_n_47));
 assign in1_85_8_ = ~((sub_781_2_n_113 & ~sub_781_2_n_152) | (sub_781_2_n_6 & sub_781_2_n_152));
 assign sub_781_2_n_154 = ~(sub_781_2_n_151 | sub_781_2_n_131);
 assign sub_781_2_n_153 = ~(sub_781_2_n_74 & (sub_781_2_n_150 | sub_781_2_n_70));
 assign sub_781_2_n_152 = ~sub_781_2_n_151;
 assign sub_781_2_n_151 = ~(sub_781_2_n_31 | sub_781_2_n_134);
 assign sub_781_2_n_150 = ~(sub_781_2_n_124 | ~(sub_781_2_n_144 | sub_781_2_n_99));
 assign sub_781_2_n_149 = ~(sub_781_2_n_42 | ~(sub_781_2_n_144 | sub_781_2_n_73));
 assign in1_85_3_ = (sub_781_2_n_145 ^ sub_781_2_n_15);
 assign sub_781_2_n_147 = ~(sub_781_2_n_146 | sub_781_2_n_141);
 assign sub_781_2_n_146 = (sub_781_2_n_143 & sub_781_2_n_129);
 assign sub_781_2_n_145 = ~(sub_781_2_n_63 & (sub_781_2_n_140 | sub_781_2_n_62));
 assign sub_781_2_n_144 = ~(sub_781_2_n_142 | sub_781_2_n_118);
 assign sub_781_2_n_143 = ~(sub_781_2_n_136 & (sub_781_2_n_135 | sub_781_2_n_123));
 assign sub_781_2_n_142 = ~(sub_781_2_n_140 | sub_781_2_n_89);
 assign sub_781_2_n_141 = ~(sub_781_2_n_133 & ~(sub_781_2_n_137 & sub_781_2_n_127));
 assign sub_781_2_n_140 = ~(sub_781_2_n_139 | sub_781_2_n_37);
 assign sub_781_2_n_139 = ~(sub_781_2_n_132 & ~(sub_781_2_n_38 & in1_83_0_));
 assign in1_85_1_ = ~(in1_83_0_ ^ (n_1586 ^ sub_781_2_n_38));
 assign sub_781_2_n_137 = ~(sub_781_2_n_115 & (sub_781_2_n_120 | sub_781_2_n_103));
 assign sub_781_2_n_136 = ~(sub_781_2_n_114 | (sub_781_2_n_125 & sub_781_2_n_108));
 assign sub_781_2_n_135 = ~(sub_781_2_n_130 | sub_781_2_n_122);
 assign sub_781_2_n_134 = ~(sub_781_2_n_116 & ~(sub_781_2_n_124 & sub_781_2_n_109));
 assign sub_781_2_n_133 = ~(sub_781_2_n_18 | sub_781_2_n_117);
 assign sub_781_2_n_132 = ~(sub_781_2_n_38 & ~n_1586);
 assign sub_781_2_n_131 = (sub_781_2_n_21 | sub_781_2_n_123);
 assign sub_781_2_n_130 = ~(sub_781_2_n_121 | sub_781_2_n_95);
 assign sub_781_2_n_129 = ~(sub_781_2_n_128 | sub_781_2_n_126);
 assign sub_781_2_n_127 = ~sub_781_2_n_126;
 assign sub_781_2_n_122 = ~(sub_781_2_n_81 & (sub_781_2_n_71 | sub_781_2_n_43));
 assign sub_781_2_n_128 = ~(sub_781_2_n_110 & sub_781_2_n_102);
 assign sub_781_2_n_126 = ~(sub_781_2_n_92 & ~sub_781_2_n_96);
 assign sub_781_2_n_125 = ~(sub_781_2_n_82 & (sub_781_2_n_76 | sub_781_2_n_44));
 assign sub_781_2_n_124 = ~(sub_781_2_n_59 & (sub_781_2_n_41 | sub_781_2_n_69));
 assign sub_781_2_n_123 = ~(sub_781_2_n_101 & sub_781_2_n_108);
 assign sub_781_2_n_118 = ~(sub_781_2_n_84 & (sub_781_2_n_63 | sub_781_2_n_49));
 assign sub_781_2_n_117 = ~(sub_781_2_n_61 & (sub_781_2_n_45 | sub_781_2_n_2));
 assign sub_781_2_n_116 = ~(sub_781_2_n_80 | ~(sub_781_2_n_74 | sub_781_2_n_64));
 assign sub_781_2_n_115 = ~(sub_781_2_n_79 | (sub_781_2_n_40 & sub_781_2_n_65));
 assign sub_781_2_n_114 = ~(sub_781_2_n_83 & (sub_781_2_n_51 | sub_781_2_n_3));
 assign sub_781_2_n_121 = ~(sub_781_2_n_58 | ~(sub_781_2_n_39 | sub_781_2_n_68));
 assign sub_781_2_n_120 = ~(sub_781_2_n_85 | ~(sub_781_2_n_78 | sub_781_2_n_1));
 assign sub_781_2_n_119 = ~(sub_781_2_n_60 | ~(sub_781_2_n_67 | sub_781_2_n_53));
 assign sub_781_2_n_113 = ~sub_781_2_n_6;
 assign sub_781_2_n_111 = ~sub_781_2_n_110;
 assign sub_781_2_n_107 = ~sub_781_2_n_106;
 assign sub_781_2_n_103 = ~sub_781_2_n_102;
 assign sub_781_2_n_112 = ~(sub_781_2_n_80 | sub_781_2_n_64);
 assign sub_781_2_n_110 = ~(sub_781_2_n_52 | sub_781_2_n_1);
 assign sub_781_2_n_109 = ~(sub_781_2_n_70 | sub_781_2_n_64);
 assign sub_781_2_n_108 = ~(sub_781_2_n_66 | sub_781_2_n_3);
 assign sub_781_2_n_106 = ~(sub_781_2_n_47 | sub_781_2_n_68);
 assign sub_781_2_n_105 = ~(sub_781_2_n_46 | sub_781_2_n_5);
 assign sub_781_2_n_104 = ~(sub_781_2_n_60 | sub_781_2_n_53);
 assign sub_781_2_n_102 = ~(sub_781_2_n_56 | sub_781_2_n_0);
 assign sub_781_2_n_101 = ~(sub_781_2_n_54 | sub_781_2_n_44);
 assign sub_781_2_n_100 = ~(sub_781_2_n_79 | sub_781_2_n_0);
 assign sub_781_2_n_99 = (sub_781_2_n_73 | sub_781_2_n_69);
 assign sub_781_2_n_89 = ~(sub_781_2_n_50 & ~sub_781_2_n_62);
 assign in1_85_0_ = ~(sub_781_2_n_38 & ~(sub_781_2_n_35 & n_1561));
 assign sub_781_2_n_98 = ~(sub_781_2_n_42 | sub_781_2_n_73);
 assign sub_781_2_n_97 = ~(sub_781_2_n_85 | sub_781_2_n_1);
 assign sub_781_2_n_96 = (sub_781_2_n_75 | sub_781_2_n_53);
 assign sub_781_2_n_95 = ~(sub_781_2_n_4 & ~sub_781_2_n_43);
 assign sub_781_2_n_94 = ~(sub_781_2_n_58 | sub_781_2_n_68);
 assign sub_781_2_n_93 = ~(sub_781_2_n_3 | ~sub_781_2_n_83);
 assign sub_781_2_n_92 = ~(sub_781_2_n_5 | sub_781_2_n_2);
 assign sub_781_2_n_87 = ~(sub_781_2_n_51 & ~sub_781_2_n_66);
 assign sub_781_2_n_91 = ~(sub_781_2_n_77 | sub_781_2_n_54);
 assign sub_781_2_n_86 = ~(sub_781_2_n_81 & ~sub_781_2_n_43);
 assign sub_781_2_n_90 = ~(sub_781_2_n_40 | sub_781_2_n_56);
 assign sub_781_2_n_77 = ~sub_781_2_n_76;
 assign sub_781_2_n_72 = ~sub_781_2_n_71;
 assign sub_781_2_n_65 = ~sub_781_2_n_0;
 assign sub_781_2_n_85 = ~(n_1562 | ~in1_83_16_);
 assign sub_781_2_n_84 = ~(in1_83_2_ & ~n_1579);
 assign sub_781_2_n_83 = ~(in1_83_14_ & ~n_1495);
 assign sub_781_2_n_82 = ~(in1_83_12_ & ~n_1581);
 assign sub_781_2_n_81 = ~(in1_83_10_ & ~n_1555);
 assign sub_781_2_n_80 = ~(n_1527 | ~in1_83_6_);
 assign sub_781_2_n_79 = ~(n_1558 | ~in1_83_18_);
 assign sub_781_2_n_78 = ~(in1_83_15_ & ~n_1549);
 assign sub_781_2_n_76 = ~(in1_83_11_ & ~n_1595);
 assign sub_781_2_n_75 = ~(in1_83_19_ | ~n_1565);
 assign sub_781_2_n_74 = ~(in1_83_5_ & ~n_1567);
 assign sub_781_2_n_73 = ~(in1_83_3_ | ~n_1535);
 assign sub_781_2_n_71 = ~(in1_83_9_ & ~n_1551);
 assign sub_781_2_n_70 = ~(in1_83_5_ | ~n_1567);
 assign sub_781_2_n_69 = ~(in1_83_4_ | ~n_1569);
 assign sub_781_2_n_68 = ~(in1_83_8_ | ~n_1589);
 assign sub_781_2_n_67 = ~(in1_83_19_ & ~n_1565);
 assign sub_781_2_n_66 = ~(in1_83_13_ | ~n_1577);
 assign sub_781_2_n_64 = ~(in1_83_6_ | ~n_1527);
 assign sub_781_2_n_63 = ~(in1_83_1_ & ~n_1477);
 assign sub_781_2_n_62 = ~(in1_83_1_ | ~n_1477);
 assign sub_781_2_n_57 = ~sub_781_2_n_56;
 assign sub_781_2_n_55 = ~sub_781_2_n_54;
 assign sub_781_2_n_50 = ~sub_781_2_n_49;
 assign sub_781_2_n_48 = ~sub_781_2_n_5;
 assign sub_781_2_n_46 = ~sub_781_2_n_45;
 assign sub_781_2_n_42 = ~sub_781_2_n_41;
 assign sub_781_2_n_37 = ~(n_1586 | ~in1_83_0_);
 assign sub_781_2_n_61 = ~(in1_83_22_ & ~n_1403);
 assign sub_781_2_n_60 = ~(n_1593 | ~in1_83_20_);
 assign sub_781_2_n_59 = ~(in1_83_4_ & ~n_1569);
 assign sub_781_2_n_58 = ~(n_1589 | ~in1_83_8_);
 assign sub_781_2_n_56 = ~(in1_83_17_ | ~n_1472);
 assign sub_781_2_n_54 = ~(in1_83_11_ | ~n_1595);
 assign sub_781_2_n_53 = ~(in1_83_20_ | ~n_1593);
 assign sub_781_2_n_52 = ~(in1_83_15_ | ~n_1549);
 assign sub_781_2_n_51 = ~(in1_83_13_ & ~n_1577);
 assign sub_781_2_n_49 = ~(in1_83_2_ | ~n_1579);
 assign sub_781_2_n_47 = ~(in1_83_7_ | ~n_1479);
 assign sub_781_2_n_45 = ~(in1_83_21_ & ~n_1591);
 assign sub_781_2_n_44 = ~(in1_83_12_ | ~n_1581);
 assign sub_781_2_n_43 = ~(in1_83_10_ | ~n_1555);
 assign sub_781_2_n_41 = ~(in1_83_3_ & ~n_1535);
 assign sub_781_2_n_40 = ~(n_1472 | ~in1_83_17_);
 assign sub_781_2_n_39 = ~(in1_83_7_ & ~n_1479);
 assign sub_781_2_n_38 = ~(n_1543 & ~n_1561);
 assign sub_781_2_n_36 = ~in1_83_23_;
 assign sub_781_2_n_35 = ~n_1543;
 assign in1_85_20_ = ~(sub_781_2_n_169 ^ sub_781_2_n_12);
 assign in1_85_7_ = (sub_781_2_n_153 ^ sub_781_2_n_112);
 assign in1_85_5_ = ~(sub_781_2_n_149 ^ sub_781_2_n_9);
 assign sub_781_2_n_31 = ~(sub_781_2_n_144 | (sub_781_2_n_99 | ~sub_781_2_n_109));
 assign in1_85_6_ = ~(sub_781_2_n_150 ^ sub_781_2_n_13);
 assign in1_85_23_ = ~(sub_781_2_n_178 ^ sub_781_2_n_10);
 assign in1_85_22_ = (sub_781_2_n_177 ^ sub_781_2_n_105);
 assign in1_85_21_ = (sub_781_2_n_176 ^ sub_781_2_n_104);
 assign in1_85_2_ = ~(sub_781_2_n_140 ^ sub_781_2_n_11);
 assign in1_85_19_ = ~(sub_781_2_n_175 ^ sub_781_2_n_100);
 assign in1_85_4_ = ~(sub_781_2_n_144 ^ sub_781_2_n_98);
 assign in1_85_17_ = (sub_781_2_n_167 ^ sub_781_2_n_97);
 assign in1_85_10_ = (sub_781_2_n_157 ^ sub_781_2_n_8);
 assign sub_781_2_n_21 = ~(sub_781_2_n_106 & ~sub_781_2_n_95);
 assign in1_85_9_ = (sub_781_2_n_156 ^ sub_781_2_n_94);
 assign in1_85_15_ = (sub_781_2_n_174 ^ sub_781_2_n_93);
 assign sub_781_2_n_18 = ~(sub_781_2_n_119 | ~sub_781_2_n_92);
 assign in1_85_12_ = (sub_781_2_n_158 ^ sub_781_2_n_91);
 assign in1_85_18_ = (sub_781_2_n_168 ^ sub_781_2_n_90);
 assign sub_781_2_n_15 = ~(sub_781_2_n_49 | ~sub_781_2_n_84);
 assign sub_781_2_n_14 = ~(sub_781_2_n_52 | ~sub_781_2_n_78);
 assign sub_781_2_n_13 = ~(sub_781_2_n_70 | ~sub_781_2_n_74);
 assign sub_781_2_n_12 = ~(sub_781_2_n_75 | ~sub_781_2_n_67);
 assign sub_781_2_n_11 = ~(sub_781_2_n_62 | ~sub_781_2_n_63);
 assign sub_781_2_n_10 = ~(sub_781_2_n_2 | ~sub_781_2_n_61);
 assign sub_781_2_n_9 = ~(sub_781_2_n_69 | ~sub_781_2_n_59);
 assign sub_781_2_n_8 = ~(sub_781_2_n_72 | ~sub_781_2_n_4);
 assign sub_781_2_n_7 = ~(sub_781_2_n_82 & ~sub_781_2_n_44);
 assign sub_781_2_n_6 = ~(sub_781_2_n_47 | ~sub_781_2_n_39);
 assign sub_781_2_n_5 = ~(in1_83_21_ | ~n_1591);
 assign sub_781_2_n_4 = ~(n_1551 & ~in1_83_9_);
 assign sub_781_2_n_3 = ~(in1_83_14_ | ~n_1495);
 assign sub_781_2_n_2 = ~(in1_83_22_ | ~n_1403);
 assign sub_781_2_n_1 = ~(in1_83_16_ | ~n_1562);
 assign sub_781_2_n_0 = ~(in1_83_18_ | ~n_1558);
 assign in1_88_23_ = ~(sub_802_2_n_182 ^ sub_802_2_n_4);
 assign sub_802_2_n_182 = ~(sub_802_2_n_178 | sub_802_2_n_43);
 assign in1_88_22_ = ~(sub_802_2_n_177 ^ sub_802_2_n_94);
 assign in1_88_19_ = ~(sub_802_2_n_174 ^ sub_802_2_n_92);
 assign in1_88_15_ = ~(sub_802_2_n_173 ^ sub_802_2_n_5);
 assign sub_802_2_n_178 = ~(sub_802_2_n_177 | sub_802_2_n_44);
 assign in1_88_24_ = ~(sub_802_2_n_162 ^ in1_86_23_);
 assign sub_802_2_n_175 = ~(sub_802_2_n_166 | sub_802_2_n_66);
 assign sub_802_2_n_174 = ~(sub_802_2_n_32 | ~(sub_802_2_n_164 | sub_802_2_n_31));
 assign sub_802_2_n_173 = ~(sub_802_2_n_165 | sub_802_2_n_34);
 assign sub_802_2_n_177 = ~(sub_802_2_n_109 | ~(sub_802_2_n_163 | sub_802_2_n_89));
 assign in1_88_20_ = ~(sub_802_2_n_163 ^ sub_802_2_n_93);
 assign in1_88_18_ = ~(sub_802_2_n_164 ^ sub_802_2_n_85);
 assign in1_88_17_ = ~(sub_802_2_n_161 ^ sub_802_2_n_3);
 assign in1_88_14_ = ~(sub_802_2_n_15 ^ sub_802_2_n_80);
 assign in1_88_13_ = ~(sub_802_2_n_156 ^ sub_802_2_n_79);
 assign in1_88_11_ = ~(sub_802_2_n_155 ^ sub_802_2_n_81);
 assign sub_802_2_n_166 = ~(sub_802_2_n_163 | sub_802_2_n_60);
 assign sub_802_2_n_165 = ~(sub_802_2_n_15 | sub_802_2_n_39);
 assign sub_802_2_n_162 = ~(sub_802_2_n_150 & sub_802_2_n_136);
 assign sub_802_2_n_161 = ~(sub_802_2_n_30 | ~(sub_802_2_n_149 | sub_802_2_n_63));
 assign sub_802_2_n_164 = ~(sub_802_2_n_14 | sub_802_2_n_110);
 assign sub_802_2_n_163 = ~(sub_802_2_n_154 | sub_802_2_n_125);
 assign in1_88_10_ = ~(sub_802_2_n_147 ^ sub_802_2_n_77);
 assign in1_88_12_ = ~(sub_802_2_n_148 ^ sub_802_2_n_82);
 assign in1_88_16_ = ~(sub_802_2_n_149 ^ sub_802_2_n_83);
 assign in1_88_9_ = ~(sub_802_2_n_146 ^ sub_802_2_n_7);
 assign sub_802_2_n_156 = ~(sub_802_2_n_152 | sub_802_2_n_38);
 assign sub_802_2_n_155 = ~(sub_802_2_n_151 | sub_802_2_n_55);
 assign sub_802_2_n_154 = ~(sub_802_2_n_149 | sub_802_2_n_115);
 assign sub_802_2_n_153 = ~(sub_802_2_n_148 | sub_802_2_n_6);
 assign sub_802_2_n_152 = ~(sub_802_2_n_148 | sub_802_2_n_52);
 assign sub_802_2_n_151 = ~(sub_802_2_n_147 | sub_802_2_n_58);
 assign sub_802_2_n_150 = ~(sub_802_2_n_131 | (sub_802_2_n_144 & sub_802_2_n_17));
 assign sub_802_2_n_149 = ~(sub_802_2_n_144 | sub_802_2_n_133);
 assign sub_802_2_n_148 = ~(sub_802_2_n_16 | sub_802_2_n_124);
 assign sub_802_2_n_147 = ~(sub_802_2_n_117 | ~(sub_802_2_n_142 | sub_802_2_n_91));
 assign sub_802_2_n_146 = ~(sub_802_2_n_70 | ~(sub_802_2_n_142 | sub_802_2_n_36));
 assign in1_88_8_ = ~(sub_802_2_n_142 ^ sub_802_2_n_78);
 assign sub_802_2_n_144 = ~(sub_802_2_n_142 | sub_802_2_n_120);
 assign sub_802_2_n_143 = ~(sub_802_2_n_54 | (sub_802_2_n_140 & sub_802_2_n_0));
 assign sub_802_2_n_142 = ~(sub_802_2_n_141 | sub_802_2_n_123);
 assign sub_802_2_n_141 = ~(sub_802_2_n_137 | sub_802_2_n_90);
 assign sub_802_2_n_140 = ~(sub_802_2_n_137 & sub_802_2_n_112);
 assign sub_802_2_n_139 = ~(sub_802_2_n_23 | (sub_802_2_n_134 & sub_802_2_n_27));
 assign in1_88_4_ = ~(sub_802_2_n_134 ^ sub_802_2_n_84);
 assign sub_802_2_n_137 = ~(sub_802_2_n_134 & sub_802_2_n_95);
 assign sub_802_2_n_136 = ~(sub_802_2_n_133 & sub_802_2_n_17);
 assign sub_802_2_n_135 = ~(sub_802_2_n_41 | (sub_802_2_n_130 & sub_802_2_n_57));
 assign sub_802_2_n_134 = ~(sub_802_2_n_132 & sub_802_2_n_114);
 assign sub_802_2_n_133 = ~(sub_802_2_n_127 & ~(sub_802_2_n_124 & sub_802_2_n_119));
 assign sub_802_2_n_132 = ~(sub_802_2_n_130 & sub_802_2_n_96);
 assign sub_802_2_n_131 = ~(sub_802_2_n_126 & ~(sub_802_2_n_125 & sub_802_2_n_118));
 assign sub_802_2_n_130 = ~(sub_802_2_n_129 & sub_802_2_n_21);
 assign sub_802_2_n_129 = ~(sub_802_2_n_122 | (sub_802_2_n_50 & in1_86_0_));
 assign in1_88_1_ = ~(in1_86_0_ ^ (n_1586 ^ sub_802_2_n_50));
 assign sub_802_2_n_127 = ~(sub_802_2_n_121 | sub_802_2_n_105);
 assign sub_802_2_n_126 = ~(sub_802_2_n_107 | (sub_802_2_n_109 & sub_802_2_n_99));
 assign sub_802_2_n_125 = ~(sub_802_2_n_108 & ~(sub_802_2_n_110 & sub_802_2_n_97));
 assign sub_802_2_n_124 = ~(sub_802_2_n_113 & ~(sub_802_2_n_117 & sub_802_2_n_100));
 assign sub_802_2_n_123 = ~(sub_802_2_n_106 & (sub_802_2_n_112 | sub_802_2_n_90));
 assign sub_802_2_n_122 = ~(n_1586 | ~sub_802_2_n_50);
 assign sub_802_2_n_121 = ~(sub_802_2_n_111 | sub_802_2_n_88);
 assign sub_802_2_n_120 = ~(sub_802_2_n_116 & sub_802_2_n_119);
 assign sub_802_2_n_114 = ~(sub_802_2_n_87 | sub_802_2_n_72);
 assign sub_802_2_n_113 = ~(sub_802_2_n_75 | (sub_802_2_n_55 & sub_802_2_n_25));
 assign sub_802_2_n_119 = ~(sub_802_2_n_6 | sub_802_2_n_88);
 assign sub_802_2_n_118 = ~(sub_802_2_n_89 | ~sub_802_2_n_99);
 assign sub_802_2_n_117 = ~(sub_802_2_n_71 & (sub_802_2_n_69 | sub_802_2_n_51));
 assign sub_802_2_n_116 = ~(sub_802_2_n_91 | ~sub_802_2_n_100);
 assign sub_802_2_n_115 = ~(sub_802_2_n_104 & sub_802_2_n_97);
 assign sub_802_2_n_108 = ~(sub_802_2_n_49 | (sub_802_2_n_32 & sub_802_2_n_67));
 assign sub_802_2_n_107 = ~(sub_802_2_n_46 & (sub_802_2_n_42 | sub_802_2_n_59));
 assign sub_802_2_n_106 = ~(sub_802_2_n_73 | ~(sub_802_2_n_53 | sub_802_2_n_28));
 assign sub_802_2_n_105 = ~(sub_802_2_n_47 & ~(sub_802_2_n_34 & sub_802_2_n_62));
 assign sub_802_2_n_112 = ~(sub_802_2_n_48 | ~(sub_802_2_n_22 | sub_802_2_n_61));
 assign sub_802_2_n_111 = ~(sub_802_2_n_76 | ~(sub_802_2_n_37 | sub_802_2_n_64));
 assign sub_802_2_n_110 = ~(sub_802_2_n_45 & (sub_802_2_n_29 | sub_802_2_n_35));
 assign sub_802_2_n_109 = ~(sub_802_2_n_74 & (sub_802_2_n_65 | sub_802_2_n_33));
 assign sub_802_2_n_96 = ~(sub_802_2_n_56 | sub_802_2_n_1);
 assign sub_802_2_n_95 = ~(sub_802_2_n_26 | sub_802_2_n_61);
 assign sub_802_2_n_104 = ~(sub_802_2_n_63 | sub_802_2_n_35);
 assign sub_802_2_n_103 = ~(sub_802_2_n_72 | sub_802_2_n_1);
 assign sub_802_2_n_102 = ~(sub_802_2_n_48 | sub_802_2_n_61);
 assign sub_802_2_n_101 = ~(sub_802_2_n_41 | sub_802_2_n_56);
 assign sub_802_2_n_100 = ~(sub_802_2_n_58 | sub_802_2_n_24);
 assign sub_802_2_n_99 = ~(sub_802_2_n_44 | sub_802_2_n_59);
 assign sub_802_2_n_94 = ~(sub_802_2_n_43 | sub_802_2_n_44);
 assign sub_802_2_n_98 = ~(sub_802_2_n_73 | sub_802_2_n_28);
 assign sub_802_2_n_97 = ~(sub_802_2_n_31 | sub_802_2_n_68);
 assign sub_802_2_n_93 = ~(sub_802_2_n_66 | sub_802_2_n_60);
 assign sub_802_2_n_92 = ~(sub_802_2_n_49 | sub_802_2_n_68);
 assign sub_802_2_n_87 = ~(sub_802_2_n_40 | sub_802_2_n_1);
 assign in1_88_0_ = ~(sub_802_2_n_50 & ~(sub_802_2_n_20 & n_1584));
 assign sub_802_2_n_85 = ~(sub_802_2_n_32 | sub_802_2_n_31);
 assign sub_802_2_n_84 = ~(sub_802_2_n_22 & sub_802_2_n_27);
 assign sub_802_2_n_83 = ~(sub_802_2_n_30 | sub_802_2_n_63);
 assign sub_802_2_n_82 = ~(sub_802_2_n_38 | sub_802_2_n_52);
 assign sub_802_2_n_81 = ~(sub_802_2_n_75 | sub_802_2_n_24);
 assign sub_802_2_n_80 = ~(sub_802_2_n_34 | sub_802_2_n_39);
 assign sub_802_2_n_91 = (sub_802_2_n_36 | sub_802_2_n_51);
 assign sub_802_2_n_79 = ~(sub_802_2_n_76 | sub_802_2_n_64);
 assign sub_802_2_n_90 = ~(sub_802_2_n_0 & ~sub_802_2_n_28);
 assign sub_802_2_n_78 = ~(sub_802_2_n_70 | sub_802_2_n_36);
 assign sub_802_2_n_77 = ~(sub_802_2_n_55 | sub_802_2_n_58);
 assign sub_802_2_n_89 = (sub_802_2_n_60 | sub_802_2_n_33);
 assign sub_802_2_n_88 = ~(sub_802_2_n_62 & ~sub_802_2_n_39);
 assign sub_802_2_n_70 = ~sub_802_2_n_69;
 assign sub_802_2_n_67 = ~sub_802_2_n_68;
 assign sub_802_2_n_66 = ~sub_802_2_n_65;
 assign sub_802_2_n_57 = ~sub_802_2_n_56;
 assign sub_802_2_n_54 = ~sub_802_2_n_53;
 assign sub_802_2_n_76 = ~(n_1581 | ~in1_86_12_);
 assign sub_802_2_n_75 = ~(n_1555 | ~in1_86_10_);
 assign sub_802_2_n_74 = ~(in1_86_20_ & ~n_1593);
 assign sub_802_2_n_73 = ~(n_1527 | ~in1_86_6_);
 assign sub_802_2_n_72 = ~(n_1579 | ~in1_86_2_);
 assign sub_802_2_n_71 = ~(in1_86_8_ & ~n_1589);
 assign sub_802_2_n_69 = ~(in1_86_7_ & ~n_1479);
 assign sub_802_2_n_68 = ~(in1_86_18_ | ~n_1558);
 assign sub_802_2_n_65 = ~(in1_86_19_ & ~n_1565);
 assign sub_802_2_n_64 = ~(in1_86_12_ | ~n_1581);
 assign sub_802_2_n_63 = ~(in1_86_15_ | ~n_1549);
 assign sub_802_2_n_62 = ~(n_1495 & ~in1_86_14_);
 assign sub_802_2_n_61 = ~(in1_86_4_ | sub_802_2_n_19);
 assign sub_802_2_n_60 = ~(in1_86_19_ | ~n_1565);
 assign sub_802_2_n_59 = ~(in1_86_22_ | ~n_1403);
 assign sub_802_2_n_58 = ~(in1_86_9_ | ~n_1551);
 assign sub_802_2_n_56 = ~(in1_86_1_ | ~n_1477);
 assign sub_802_2_n_55 = ~(n_1551 | ~in1_86_9_);
 assign sub_802_2_n_53 = ~(in1_86_5_ & ~n_1567);
 assign sub_802_2_n_52 = ~(in1_86_11_ | ~n_1595);
 assign sub_802_2_n_51 = ~(in1_86_8_ | ~n_1589);
 assign sub_802_2_n_50 = ~(n_1543 & ~n_1584);
 assign sub_802_2_n_43 = ~sub_802_2_n_42;
 assign sub_802_2_n_41 = ~sub_802_2_n_40;
 assign sub_802_2_n_38 = ~sub_802_2_n_37;
 assign sub_802_2_n_30 = ~sub_802_2_n_29;
 assign sub_802_2_n_27 = ~sub_802_2_n_26;
 assign sub_802_2_n_25 = ~sub_802_2_n_24;
 assign sub_802_2_n_23 = ~sub_802_2_n_22;
 assign sub_802_2_n_21 = ~(in1_86_0_ & ~n_1586);
 assign sub_802_2_n_49 = ~(n_1558 | ~in1_86_18_);
 assign sub_802_2_n_48 = (sub_802_2_n_19 & in1_86_4_);
 assign sub_802_2_n_47 = ~(in1_86_14_ & ~n_1495);
 assign sub_802_2_n_46 = ~(in1_86_22_ & ~n_1403);
 assign sub_802_2_n_45 = ~(in1_86_16_ & ~n_1562);
 assign sub_802_2_n_44 = ~(in1_86_21_ | ~n_1591);
 assign sub_802_2_n_42 = ~(in1_86_21_ & ~n_1591);
 assign sub_802_2_n_40 = ~(in1_86_1_ & ~n_1477);
 assign sub_802_2_n_39 = ~(in1_86_13_ | ~n_1577);
 assign sub_802_2_n_37 = ~(in1_86_11_ & ~n_1595);
 assign sub_802_2_n_36 = ~(in1_86_7_ | ~n_1479);
 assign sub_802_2_n_35 = ~(in1_86_16_ | ~n_1562);
 assign sub_802_2_n_34 = ~(n_1577 | ~in1_86_13_);
 assign sub_802_2_n_33 = ~(in1_86_20_ | ~n_1593);
 assign sub_802_2_n_32 = ~(n_1472 | ~in1_86_17_);
 assign sub_802_2_n_31 = ~(in1_86_17_ | ~n_1472);
 assign sub_802_2_n_29 = ~(in1_86_15_ & ~n_1549);
 assign sub_802_2_n_28 = ~(in1_86_6_ | ~n_1527);
 assign sub_802_2_n_26 = ~(in1_86_3_ | ~n_1535);
 assign sub_802_2_n_24 = ~(in1_86_10_ | ~n_1555);
 assign sub_802_2_n_22 = ~(in1_86_3_ & ~n_1535);
 assign sub_802_2_n_20 = ~n_1543;
 assign sub_802_2_n_19 = ~n_1569;
 assign in1_88_6_ = (sub_802_2_n_140 ^ sub_802_2_n_2);
 assign sub_802_2_n_17 = ~(sub_802_2_n_115 | ~sub_802_2_n_118);
 assign sub_802_2_n_16 = ~(sub_802_2_n_142 | ~sub_802_2_n_116);
 assign sub_802_2_n_15 = ~(sub_802_2_n_153 | ~sub_802_2_n_111);
 assign sub_802_2_n_14 = ~(sub_802_2_n_149 | ~sub_802_2_n_104);
 assign in1_88_3_ = ~(sub_802_2_n_135 ^ sub_802_2_n_103);
 assign in1_88_5_ = ~(sub_802_2_n_139 ^ sub_802_2_n_102);
 assign in1_88_2_ = (sub_802_2_n_130 ^ sub_802_2_n_101);
 assign in1_88_21_ = ~(sub_802_2_n_175 ^ sub_802_2_n_8);
 assign in1_88_7_ = ~(sub_802_2_n_143 ^ sub_802_2_n_98);
 assign sub_802_2_n_8 = ~(sub_802_2_n_33 | ~sub_802_2_n_74);
 assign sub_802_2_n_7 = ~(sub_802_2_n_51 | ~sub_802_2_n_71);
 assign sub_802_2_n_6 = (sub_802_2_n_64 | sub_802_2_n_52);
 assign sub_802_2_n_5 = (sub_802_2_n_47 & sub_802_2_n_62);
 assign sub_802_2_n_4 = ~(sub_802_2_n_59 | ~sub_802_2_n_46);
 assign sub_802_2_n_3 = ~(sub_802_2_n_35 | ~sub_802_2_n_45);
 assign sub_802_2_n_2 = ~(sub_802_2_n_54 | ~sub_802_2_n_0);
 assign sub_802_2_n_1 = ~(in1_86_2_ | ~n_1579);
 assign sub_802_2_n_0 = ~(n_1567 & ~in1_86_5_);
 assign sub_823_2_n_173 = ~(sub_823_2_n_51 & (sub_823_2_n_172 | sub_823_2_n_3));
 assign sub_823_2_n_172 = ~(sub_823_2_n_116 | (sub_823_2_n_36 & sub_823_2_n_97));
 assign sub_823_2_n_171 = ~(sub_823_2_n_73 & (sub_823_2_n_165 | sub_823_2_n_2));
 assign sub_823_2_n_170 = ~(sub_823_2_n_77 & (sub_823_2_n_164 | sub_823_2_n_53));
 assign in1_91_18_ = (sub_823_2_n_164 ^ sub_823_2_n_88);
 assign sub_823_2_n_168 = ~(sub_823_2_n_47 & (sub_823_2_n_158 | sub_823_2_n_58));
 assign in1_91_24_ = ~(sub_823_2_n_166 & (sub_823_2_n_159 | in1_89_23_));
 assign sub_823_2_n_166 = ~(sub_823_2_n_159 & in1_89_23_);
 assign sub_823_2_n_165 = ~sub_823_2_n_36;
 assign sub_823_2_n_164 = ~(sub_823_2_n_160 | sub_823_2_n_117);
 assign sub_823_2_n_163 = ~(sub_823_2_n_75 & (sub_823_2_n_154 | sub_823_2_n_50));
 assign in1_91_16_ = (sub_823_2_n_154 ^ sub_823_2_n_87);
 assign sub_823_2_n_161 = ~(sub_823_2_n_40 & sub_823_2_n_24);
 assign sub_823_2_n_160 = ~(sub_823_2_n_154 | sub_823_2_n_98);
 assign sub_823_2_n_159 = ~(sub_823_2_n_141 & sub_823_2_n_155);
 assign sub_823_2_n_158 = ~(sub_823_2_n_25 | sub_823_2_n_121);
 assign sub_823_2_n_157 = ~(sub_823_2_n_76 & (sub_823_2_n_39 | sub_823_2_n_54));
 assign in1_91_12_ = ~(sub_823_2_n_39 ^ sub_823_2_n_15);
 assign sub_823_2_n_155 = ~(sub_823_2_n_151 & sub_823_2_n_124);
 assign sub_823_2_n_154 = ~sub_823_2_n_40;
 assign sub_823_2_n_153 = ~(sub_823_2_n_70 & (sub_823_2_n_34 | sub_823_2_n_48));
 assign in1_91_10_ = (sub_823_2_n_34 ^ sub_823_2_n_91);
 assign sub_823_2_n_151 = ~(sub_823_2_n_20 | sub_823_2_n_120);
 assign in1_91_7_ = (sub_823_2_n_148 ^ sub_823_2_n_90);
 assign sub_823_2_n_149 = ~(sub_823_2_n_56 & (sub_823_2_n_146 | sub_823_2_n_55));
 assign sub_823_2_n_148 = ~(sub_823_2_n_72 & (sub_823_2_n_37 | sub_823_2_n_0));
 assign sub_823_2_n_147 = ~(sub_823_2_n_146 | sub_823_2_n_93);
 assign sub_823_2_n_146 = ~(sub_823_2_n_31 | sub_823_2_n_129);
 assign sub_823_2_n_145 = ~(sub_823_2_n_81 | (sub_823_2_n_138 & sub_823_2_n_68));
 assign in1_91_4_ = ~(sub_823_2_n_138 ^ sub_823_2_n_101);
 assign in1_91_3_ = (sub_823_2_n_139 ^ sub_823_2_n_89);
 assign sub_823_2_n_142 = ~(sub_823_2_n_138 & sub_823_2_n_102);
 assign sub_823_2_n_141 = ~(sub_823_2_n_140 | sub_823_2_n_135);
 assign sub_823_2_n_140 = ~(sub_823_2_n_136 | ~sub_823_2_n_124);
 assign sub_823_2_n_139 = ~(sub_823_2_n_52 & (sub_823_2_n_133 | sub_823_2_n_74));
 assign sub_823_2_n_138 = ~(sub_823_2_n_137 & sub_823_2_n_112);
 assign sub_823_2_n_137 = ~(sub_823_2_n_134 & sub_823_2_n_94);
 assign sub_823_2_n_136 = ~(sub_823_2_n_131 | sub_823_2_n_127);
 assign sub_823_2_n_135 = ~(sub_823_2_n_35 & sub_823_2_n_126);
 assign sub_823_2_n_133 = ~sub_823_2_n_134;
 assign sub_823_2_n_134 = ((sub_823_2_n_45 & in1_89_0_) | ((in1_89_0_ & sub_823_2_n_43) | (sub_823_2_n_43
    & sub_823_2_n_45)));
 assign in1_91_1_ = (in1_89_0_ ^ (sub_823_2_n_43 ^ sub_823_2_n_45));
 assign sub_823_2_n_131 = ~(sub_823_2_n_128 | sub_823_2_n_120);
 assign sub_823_2_n_130 = ~(sub_823_2_n_113 & ~(sub_823_2_n_117 & sub_823_2_n_105));
 assign sub_823_2_n_129 = ~(sub_823_2_n_114 & ~(sub_823_2_n_115 & sub_823_2_n_109));
 assign sub_823_2_n_128 = ~(sub_823_2_n_125 | sub_823_2_n_118);
 assign sub_823_2_n_127 = ~(sub_823_2_n_119 & ~(sub_823_2_n_121 & sub_823_2_n_110));
 assign sub_823_2_n_126 = ~(sub_823_2_n_29 | sub_823_2_n_111);
 assign sub_823_2_n_125 = ~(sub_823_2_n_122 | sub_823_2_n_100);
 assign sub_823_2_n_124 = ~(sub_823_2_n_123 | ~sub_823_2_n_24);
 assign sub_823_2_n_119 = ~(sub_823_2_n_64 | ~(sub_823_2_n_47 | sub_823_2_n_69));
 assign sub_823_2_n_118 = ~(sub_823_2_n_82 & (sub_823_2_n_70 | sub_823_2_n_59));
 assign sub_823_2_n_123 = ~(sub_823_2_n_97 & sub_823_2_n_108);
 assign sub_823_2_n_122 = ~(sub_823_2_n_103 | sub_823_2_n_60);
 assign sub_823_2_n_121 = ~(sub_823_2_n_62 & (sub_823_2_n_76 | sub_823_2_n_49));
 assign sub_823_2_n_120 = ~(sub_823_2_n_106 & sub_823_2_n_110);
 assign sub_823_2_n_114 = ~(sub_823_2_n_83 | ~(sub_823_2_n_72 | sub_823_2_n_66));
 assign sub_823_2_n_113 = ~(sub_823_2_n_85 | ~(sub_823_2_n_77 | sub_823_2_n_57));
 assign sub_823_2_n_112 = ~(sub_823_2_n_86 | ~(sub_823_2_n_52 | sub_823_2_n_78));
 assign sub_823_2_n_111 = ~(sub_823_2_n_63 & (sub_823_2_n_51 | sub_823_2_n_1));
 assign sub_823_2_n_117 = ~(sub_823_2_n_84 & (sub_823_2_n_75 | sub_823_2_n_46));
 assign sub_823_2_n_116 = ~(sub_823_2_n_61 & (sub_823_2_n_73 | sub_823_2_n_71));
 assign sub_823_2_n_115 = ~(sub_823_2_n_65 & (sub_823_2_n_80 | sub_823_2_n_4));
 assign sub_823_2_n_103 = ~(sub_823_2_n_56 | sub_823_2_n_79);
 assign sub_823_2_n_102 = ~(sub_823_2_n_67 | sub_823_2_n_4);
 assign sub_823_2_n_110 = ~(sub_823_2_n_58 | sub_823_2_n_69);
 assign sub_823_2_n_109 = ~(sub_823_2_n_0 | sub_823_2_n_66);
 assign sub_823_2_n_108 = ~(sub_823_2_n_3 | sub_823_2_n_1);
 assign sub_823_2_n_107 = ~(sub_823_2_n_59 | ~sub_823_2_n_82);
 assign sub_823_2_n_106 = ~(sub_823_2_n_54 | sub_823_2_n_49);
 assign sub_823_2_n_105 = ~(sub_823_2_n_53 | sub_823_2_n_57);
 assign sub_823_2_n_104 = ~(sub_823_2_n_85 | sub_823_2_n_57);
 assign sub_823_2_n_101 = ~(sub_823_2_n_80 & sub_823_2_n_68);
 assign sub_823_2_n_94 = ~(sub_823_2_n_74 | sub_823_2_n_78);
 assign sub_823_2_n_93 = (sub_823_2_n_55 | sub_823_2_n_79);
 assign in1_91_0_ = ~(sub_823_2_n_45 & ~(sub_823_2_n_44 & n_1532));
 assign sub_823_2_n_91 = ~(sub_823_2_n_70 & ~sub_823_2_n_48);
 assign sub_823_2_n_100 = (sub_823_2_n_48 | sub_823_2_n_59);
 assign sub_823_2_n_90 = ~(sub_823_2_n_83 | sub_823_2_n_66);
 assign sub_823_2_n_89 = ~(sub_823_2_n_86 | sub_823_2_n_78);
 assign sub_823_2_n_99 = ~(sub_823_2_n_64 | sub_823_2_n_69);
 assign sub_823_2_n_88 = ~(sub_823_2_n_77 & ~sub_823_2_n_53);
 assign sub_823_2_n_87 = ~(sub_823_2_n_75 & ~sub_823_2_n_50);
 assign sub_823_2_n_98 = (sub_823_2_n_50 | sub_823_2_n_46);
 assign sub_823_2_n_97 = ~(sub_823_2_n_2 | sub_823_2_n_71);
 assign sub_823_2_n_96 = ~(sub_823_2_n_60 | sub_823_2_n_79);
 assign sub_823_2_n_95 = ~(sub_823_2_n_46 | ~sub_823_2_n_84);
 assign sub_823_2_n_81 = ~sub_823_2_n_80;
 assign sub_823_2_n_68 = ~sub_823_2_n_67;
 assign sub_823_2_n_86 = ~(n_1579 | ~in1_89_2_);
 assign sub_823_2_n_85 = ~(n_1558 | ~in1_89_18_);
 assign sub_823_2_n_84 = ~(in1_89_16_ & ~n_1562);
 assign sub_823_2_n_83 = ~(n_1527 | ~in1_89_6_);
 assign sub_823_2_n_82 = ~(in1_89_10_ & ~n_1555);
 assign sub_823_2_n_80 = ~(in1_89_3_ & ~n_1535);
 assign sub_823_2_n_79 = ~(in1_89_8_ | sub_823_2_n_42);
 assign sub_823_2_n_78 = ~(in1_89_2_ | ~n_1579);
 assign sub_823_2_n_77 = ~(in1_89_17_ & ~n_1472);
 assign sub_823_2_n_76 = ~(in1_89_11_ & ~n_1595);
 assign sub_823_2_n_75 = ~(in1_89_15_ & ~n_1549);
 assign sub_823_2_n_74 = ~(in1_89_1_ | ~n_1477);
 assign sub_823_2_n_73 = ~(in1_89_19_ & ~n_1565);
 assign sub_823_2_n_72 = ~(in1_89_5_ & ~n_1567);
 assign sub_823_2_n_71 = ~(in1_89_20_ | ~n_1593);
 assign sub_823_2_n_70 = ~(in1_89_9_ & ~n_1551);
 assign sub_823_2_n_69 = ~(in1_89_14_ | ~n_1495);
 assign sub_823_2_n_67 = ~(in1_89_3_ | ~n_1535);
 assign sub_823_2_n_66 = ~(in1_89_6_ | ~n_1527);
 assign sub_823_2_n_65 = ~(in1_89_4_ & ~n_1569);
 assign sub_823_2_n_64 = ~(n_1495 | ~in1_89_14_);
 assign sub_823_2_n_63 = ~(in1_89_22_ & ~n_1403);
 assign sub_823_2_n_62 = ~(in1_89_12_ & ~n_1581);
 assign sub_823_2_n_61 = ~(in1_89_20_ & ~n_1593);
 assign sub_823_2_n_60 = (sub_823_2_n_42 & in1_89_8_);
 assign sub_823_2_n_59 = ~(in1_89_10_ | ~n_1555);
 assign sub_823_2_n_58 = ~(in1_89_13_ | ~n_1577);
 assign sub_823_2_n_57 = ~(in1_89_18_ | ~n_1558);
 assign sub_823_2_n_56 = ~(in1_89_7_ & ~n_1479);
 assign sub_823_2_n_55 = ~(in1_89_7_ | ~n_1479);
 assign sub_823_2_n_54 = ~(in1_89_11_ | ~n_1595);
 assign sub_823_2_n_53 = ~(in1_89_17_ | ~n_1472);
 assign sub_823_2_n_52 = ~(in1_89_1_ & ~n_1477);
 assign sub_823_2_n_51 = ~(in1_89_21_ & ~n_1591);
 assign sub_823_2_n_50 = ~(in1_89_15_ | ~n_1549);
 assign sub_823_2_n_49 = ~(in1_89_12_ | ~n_1581);
 assign sub_823_2_n_48 = ~(in1_89_9_ | ~n_1551);
 assign sub_823_2_n_47 = ~(in1_89_13_ & ~n_1577);
 assign sub_823_2_n_46 = ~(in1_89_16_ | ~n_1562);
 assign sub_823_2_n_45 = ~(n_1543 & ~n_1532);
 assign sub_823_2_n_44 = ~n_1543;
 assign sub_823_2_n_43 = ~n_1586;
 assign sub_823_2_n_42 = ~n_1589;
 assign in1_91_14_ = ~(sub_823_2_n_158 ^ sub_823_2_n_5);
 assign sub_823_2_n_40 = ~(sub_823_2_n_136 & ~sub_823_2_n_151);
 assign sub_823_2_n_39 = (sub_823_2_n_20 & sub_823_2_n_128);
 assign in1_91_8_ = ~(sub_823_2_n_146 ^ sub_823_2_n_8);
 assign sub_823_2_n_37 = ~(sub_823_2_n_115 | ~sub_823_2_n_142);
 assign sub_823_2_n_36 = ~(sub_823_2_n_161 & ~sub_823_2_n_130);
 assign sub_823_2_n_35 = ~(sub_823_2_n_130 & ~sub_823_2_n_123);
 assign sub_823_2_n_34 = ~(sub_823_2_n_147 | ~sub_823_2_n_122);
 assign in1_91_23_ = (sub_823_2_n_173 ^ sub_823_2_n_11);
 assign in1_91_6_ = ~(sub_823_2_n_37 ^ sub_823_2_n_13);
 assign sub_823_2_n_31 = ~(sub_823_2_n_142 | ~sub_823_2_n_109);
 assign in1_91_5_ = ~(sub_823_2_n_145 ^ sub_823_2_n_12);
 assign sub_823_2_n_29 = (sub_823_2_n_108 & sub_823_2_n_116);
 assign in1_91_22_ = ~(sub_823_2_n_172 ^ sub_823_2_n_6);
 assign in1_91_21_ = (sub_823_2_n_171 ^ sub_823_2_n_9);
 assign in1_91_11_ = (sub_823_2_n_153 ^ sub_823_2_n_107);
 assign sub_823_2_n_25 = ~(sub_823_2_n_39 | ~sub_823_2_n_106);
 assign sub_823_2_n_24 = ~(sub_823_2_n_98 | ~sub_823_2_n_105);
 assign in1_91_2_ = (sub_823_2_n_134 ^ sub_823_2_n_7);
 assign in1_91_20_ = (sub_823_2_n_36 ^ sub_823_2_n_14);
 assign in1_91_19_ = (sub_823_2_n_170 ^ sub_823_2_n_104);
 assign sub_823_2_n_20 = ~(sub_823_2_n_147 & ~sub_823_2_n_100);
 assign in1_91_15_ = (sub_823_2_n_168 ^ sub_823_2_n_99);
 assign in1_91_13_ = (sub_823_2_n_157 ^ sub_823_2_n_10);
 assign in1_91_9_ = (sub_823_2_n_149 ^ sub_823_2_n_96);
 assign in1_91_17_ = (sub_823_2_n_163 ^ sub_823_2_n_95);
 assign sub_823_2_n_15 = ~(sub_823_2_n_54 | ~sub_823_2_n_76);
 assign sub_823_2_n_14 = ~(sub_823_2_n_2 | ~sub_823_2_n_73);
 assign sub_823_2_n_13 = ~(sub_823_2_n_0 | ~sub_823_2_n_72);
 assign sub_823_2_n_12 = ~(sub_823_2_n_4 | ~sub_823_2_n_65);
 assign sub_823_2_n_11 = ~(sub_823_2_n_1 | ~sub_823_2_n_63);
 assign sub_823_2_n_10 = ~(sub_823_2_n_49 | ~sub_823_2_n_62);
 assign sub_823_2_n_9 = ~(sub_823_2_n_71 | ~sub_823_2_n_61);
 assign sub_823_2_n_8 = ~(sub_823_2_n_55 | ~sub_823_2_n_56);
 assign sub_823_2_n_7 = ~(sub_823_2_n_74 | ~sub_823_2_n_52);
 assign sub_823_2_n_6 = ~(sub_823_2_n_3 | ~sub_823_2_n_51);
 assign sub_823_2_n_5 = ~(sub_823_2_n_58 | ~sub_823_2_n_47);
 assign sub_823_2_n_4 = ~(in1_89_4_ | ~n_1569);
 assign sub_823_2_n_3 = ~(in1_89_21_ | ~n_1591);
 assign sub_823_2_n_2 = ~(in1_89_19_ | ~n_1565);
 assign sub_823_2_n_1 = ~(in1_89_22_ | ~n_1403);
 assign sub_823_2_n_0 = ~(in1_89_5_ | ~n_1567);
 assign sub_844_2_n_171 = ~(sub_844_2_n_46 & (sub_844_2_n_169 | sub_844_2_n_69));
 assign in1_94_19_ = ~(sub_844_2_n_167 ^ sub_844_2_n_99);
 assign sub_844_2_n_169 = ~(sub_844_2_n_115 | (sub_844_2_n_162 & sub_844_2_n_102));
 assign sub_844_2_n_168 = ~(sub_844_2_n_45 & ~(sub_844_2_n_162 & sub_844_2_n_79));
 assign sub_844_2_n_167 = ~(sub_844_2_n_57 & (sub_844_2_n_161 | sub_844_2_n_73));
 assign sub_844_2_n_166 = ~(sub_844_2_n_82 & (sub_844_2_n_159 | sub_844_2_n_65));
 assign in1_94_20_ = ~(sub_844_2_n_162 ^ sub_844_2_n_100);
 assign in1_94_14_ = ~(sub_844_2_n_159 ^ sub_844_2_n_15);
 assign in1_94_24_ = ~(sub_844_2_n_156 ^ in1_92_23_);
 assign sub_844_2_n_162 = ~(sub_844_2_n_129 & (sub_844_2_n_153 | sub_844_2_n_121));
 assign sub_844_2_n_161 = ~(sub_844_2_n_20 | sub_844_2_n_114);
 assign sub_844_2_n_160 = ~(sub_844_2_n_58 & (sub_844_2_n_153 | sub_844_2_n_49));
 assign sub_844_2_n_159 = ~(sub_844_2_n_116 | (sub_844_2_n_152 & sub_844_2_n_104));
 assign sub_844_2_n_158 = ~(sub_844_2_n_77 & ~(sub_844_2_n_152 & sub_844_2_n_71));
 assign sub_844_2_n_157 = ~(sub_844_2_n_72 & (sub_844_2_n_151 | sub_844_2_n_2));
 assign sub_844_2_n_156 = ~(sub_844_2_n_154 & sub_844_2_n_141);
 assign in1_94_7_ = (sub_844_2_n_149 ^ sub_844_2_n_89);
 assign sub_844_2_n_154 = ~(sub_844_2_n_148 & sub_844_2_n_35);
 assign sub_844_2_n_153 = ~(sub_844_2_n_148 | sub_844_2_n_137);
 assign sub_844_2_n_152 = ~(sub_844_2_n_132 & (sub_844_2_n_147 | sub_844_2_n_123));
 assign sub_844_2_n_151 = ~(sub_844_2_n_113 | (sub_844_2_n_146 & sub_844_2_n_96));
 assign sub_844_2_n_150 = ~(sub_844_2_n_50 & (sub_844_2_n_147 | sub_844_2_n_75));
 assign sub_844_2_n_149 = ~(sub_844_2_n_74 & (sub_844_2_n_36 | sub_844_2_n_80));
 assign sub_844_2_n_148 = ~(sub_844_2_n_147 | sub_844_2_n_127);
 assign sub_844_2_n_146 = ~sub_844_2_n_147;
 assign sub_844_2_n_147 = ~(sub_844_2_n_145 | sub_844_2_n_131);
 assign sub_844_2_n_145 = ~(sub_844_2_n_142 | sub_844_2_n_13);
 assign sub_844_2_n_144 = ~(sub_844_2_n_51 | (sub_844_2_n_139 & sub_844_2_n_56));
 assign in1_94_4_ = ~(sub_844_2_n_139 ^ sub_844_2_n_5);
 assign sub_844_2_n_142 = ~(sub_844_2_n_139 & sub_844_2_n_101);
 assign sub_844_2_n_141 = ~(sub_844_2_n_136 | (sub_844_2_n_137 & sub_844_2_n_35));
 assign sub_844_2_n_140 = ~(sub_844_2_n_43 | (sub_844_2_n_135 & sub_844_2_n_48));
 assign sub_844_2_n_139 = ~(sub_844_2_n_138 & sub_844_2_n_110);
 assign sub_844_2_n_138 = ~(sub_844_2_n_135 & sub_844_2_n_91);
 assign sub_844_2_n_137 = ~(sub_844_2_n_130 & (sub_844_2_n_132 | sub_844_2_n_124));
 assign sub_844_2_n_136 = ~(sub_844_2_n_133 & sub_844_2_n_128);
 assign sub_844_2_n_135 = ((sub_844_2_n_41 & in1_92_0_) | ((in1_92_0_ & sub_844_2_n_40) | (sub_844_2_n_40
    & sub_844_2_n_41)));
 assign in1_94_1_ = (in1_92_0_ ^ (sub_844_2_n_40 ^ sub_844_2_n_41));
 assign sub_844_2_n_133 = ~(sub_844_2_n_122 & ~sub_844_2_n_129);
 assign sub_844_2_n_132 = ~(sub_844_2_n_24 | sub_844_2_n_111);
 assign sub_844_2_n_131 = ~(sub_844_2_n_126 & sub_844_2_n_119);
 assign sub_844_2_n_130 = ~(sub_844_2_n_120 | (sub_844_2_n_116 & sub_844_2_n_107));
 assign sub_844_2_n_129 = ~(sub_844_2_n_118 | (sub_844_2_n_114 & sub_844_2_n_105));
 assign sub_844_2_n_128 = ~(sub_844_2_n_125 | sub_844_2_n_109);
 assign sub_844_2_n_127 = (sub_844_2_n_123 | sub_844_2_n_124);
 assign sub_844_2_n_126 = ~(sub_844_2_n_117 & ~sub_844_2_n_13);
 assign sub_844_2_n_125 = ~(sub_844_2_n_106 | ~sub_844_2_n_115);
 assign sub_844_2_n_120 = ~(sub_844_2_n_62 & (sub_844_2_n_82 | sub_844_2_n_54));
 assign sub_844_2_n_119 = ~(sub_844_2_n_64 | ~(sub_844_2_n_74 | sub_844_2_n_76));
 assign sub_844_2_n_118 = ~(sub_844_2_n_87 & (sub_844_2_n_57 | sub_844_2_n_44));
 assign sub_844_2_n_124 = ~(sub_844_2_n_104 & sub_844_2_n_107);
 assign sub_844_2_n_123 = ~(sub_844_2_n_96 & sub_844_2_n_97);
 assign sub_844_2_n_122 = ~(sub_844_2_n_106 | ~sub_844_2_n_102);
 assign sub_844_2_n_121 = ~(sub_844_2_n_94 & sub_844_2_n_105);
 assign sub_844_2_n_113 = ~sub_844_2_n_112;
 assign sub_844_2_n_111 = ~(sub_844_2_n_86 & (sub_844_2_n_72 | sub_844_2_n_0));
 assign sub_844_2_n_110 = ~(sub_844_2_n_92 | sub_844_2_n_88);
 assign sub_844_2_n_109 = ~(sub_844_2_n_61 & (sub_844_2_n_46 | sub_844_2_n_81));
 assign sub_844_2_n_117 = ~(sub_844_2_n_60 & ~(sub_844_2_n_51 & sub_844_2_n_52));
 assign sub_844_2_n_116 = ~(sub_844_2_n_85 & (sub_844_2_n_77 | sub_844_2_n_59));
 assign sub_844_2_n_115 = ~(sub_844_2_n_63 & (sub_844_2_n_45 | sub_844_2_n_66));
 assign sub_844_2_n_114 = ~(sub_844_2_n_83 & (sub_844_2_n_58 | sub_844_2_n_67));
 assign sub_844_2_n_112 = ~(sub_844_2_n_84 | ~(sub_844_2_n_50 | sub_844_2_n_68));
 assign sub_844_2_n_101 = ~(sub_844_2_n_55 | sub_844_2_n_53);
 assign sub_844_2_n_108 = ~(sub_844_2_n_84 | sub_844_2_n_68);
 assign sub_844_2_n_107 = ~(sub_844_2_n_65 | sub_844_2_n_54);
 assign sub_844_2_n_106 = (sub_844_2_n_69 | sub_844_2_n_81);
 assign sub_844_2_n_105 = ~(sub_844_2_n_73 | sub_844_2_n_44);
 assign sub_844_2_n_104 = ~(sub_844_2_n_70 | sub_844_2_n_59);
 assign sub_844_2_n_100 = ~(sub_844_2_n_45 & sub_844_2_n_79);
 assign sub_844_2_n_103 = ~(sub_844_2_n_43 | sub_844_2_n_47);
 assign sub_844_2_n_99 = ~(sub_844_2_n_87 & ~sub_844_2_n_44);
 assign sub_844_2_n_102 = ~(sub_844_2_n_78 | sub_844_2_n_66);
 assign sub_844_2_n_92 = ~(sub_844_2_n_42 | sub_844_2_n_1);
 assign sub_844_2_n_91 = ~(sub_844_2_n_47 | sub_844_2_n_1);
 assign in1_94_0_ = ~(sub_844_2_n_41 & ~(sub_844_2_n_39 & n_1557));
 assign sub_844_2_n_98 = ~(sub_844_2_n_0 | ~sub_844_2_n_86);
 assign sub_844_2_n_97 = ~(sub_844_2_n_2 | sub_844_2_n_0);
 assign sub_844_2_n_96 = ~(sub_844_2_n_75 | sub_844_2_n_68);
 assign sub_844_2_n_95 = ~(sub_844_2_n_88 | sub_844_2_n_1);
 assign sub_844_2_n_89 = ~(sub_844_2_n_64 | sub_844_2_n_76);
 assign sub_844_2_n_94 = ~(sub_844_2_n_49 | sub_844_2_n_67);
 assign sub_844_2_n_93 = ~(sub_844_2_n_54 | ~sub_844_2_n_62);
 assign sub_844_2_n_79 = ~sub_844_2_n_78;
 assign sub_844_2_n_71 = ~sub_844_2_n_70;
 assign sub_844_2_n_88 = ~(n_1579 | ~in1_92_2_);
 assign sub_844_2_n_87 = ~(in1_92_18_ & ~n_1558);
 assign sub_844_2_n_86 = ~(in1_92_10_ & ~n_1555);
 assign sub_844_2_n_85 = ~(in1_92_12_ & ~n_1581);
 assign sub_844_2_n_84 = ~(n_1589 | ~in1_92_8_);
 assign sub_844_2_n_83 = ~(in1_92_16_ & ~n_1562);
 assign sub_844_2_n_82 = ~(in1_92_13_ & ~n_1577);
 assign sub_844_2_n_81 = ~(in1_92_22_ | ~n_1403);
 assign sub_844_2_n_80 = ~(in1_92_5_ | ~n_1567);
 assign sub_844_2_n_78 = ~(in1_92_19_ | ~n_1565);
 assign sub_844_2_n_77 = ~(in1_92_11_ & ~n_1595);
 assign sub_844_2_n_76 = ~(in1_92_6_ | ~n_1527);
 assign sub_844_2_n_75 = ~(in1_92_7_ | ~n_1479);
 assign sub_844_2_n_74 = ~(in1_92_5_ & ~n_1567);
 assign sub_844_2_n_73 = ~(in1_92_17_ | ~n_1472);
 assign sub_844_2_n_72 = ~(in1_92_9_ & ~n_1551);
 assign sub_844_2_n_70 = ~(in1_92_11_ | ~n_1595);
 assign sub_844_2_n_69 = ~(in1_92_21_ | ~n_1591);
 assign sub_844_2_n_68 = ~(in1_92_8_ | ~n_1589);
 assign sub_844_2_n_67 = ~(in1_92_16_ | ~n_1562);
 assign sub_844_2_n_66 = ~(in1_92_20_ | ~n_1593);
 assign sub_844_2_n_65 = ~(in1_92_13_ | ~n_1577);
 assign sub_844_2_n_56 = ~sub_844_2_n_55;
 assign sub_844_2_n_53 = ~sub_844_2_n_52;
 assign sub_844_2_n_48 = ~sub_844_2_n_47;
 assign sub_844_2_n_43 = ~sub_844_2_n_42;
 assign sub_844_2_n_64 = ~(n_1527 | ~in1_92_6_);
 assign sub_844_2_n_63 = ~(in1_92_20_ & ~n_1593);
 assign sub_844_2_n_62 = ~(in1_92_14_ & ~n_1495);
 assign sub_844_2_n_61 = ~(in1_92_22_ & ~n_1403);
 assign sub_844_2_n_60 = ~(in1_92_4_ & ~n_1569);
 assign sub_844_2_n_59 = ~(in1_92_12_ | ~n_1581);
 assign sub_844_2_n_58 = ~(in1_92_15_ & ~n_1549);
 assign sub_844_2_n_57 = ~(in1_92_17_ & ~n_1472);
 assign sub_844_2_n_55 = ~(in1_92_3_ | ~n_1535);
 assign sub_844_2_n_54 = ~(in1_92_14_ | ~n_1495);
 assign sub_844_2_n_52 = ~(n_1569 & ~in1_92_4_);
 assign sub_844_2_n_51 = ~(n_1535 | ~in1_92_3_);
 assign sub_844_2_n_50 = ~(in1_92_7_ & ~n_1479);
 assign sub_844_2_n_49 = ~(in1_92_15_ | ~n_1549);
 assign sub_844_2_n_47 = ~(in1_92_1_ | ~n_1477);
 assign sub_844_2_n_46 = ~(in1_92_21_ & ~n_1591);
 assign sub_844_2_n_45 = ~(in1_92_19_ & ~n_1565);
 assign sub_844_2_n_44 = ~(in1_92_18_ | ~n_1558);
 assign sub_844_2_n_42 = ~(in1_92_1_ & ~n_1477);
 assign sub_844_2_n_41 = ~(n_1543 & ~n_1557);
 assign sub_844_2_n_40 = ~n_1586;
 assign sub_844_2_n_39 = ~n_1543;
 assign in1_94_18_ = ~(sub_844_2_n_161 ^ sub_844_2_n_6);
 assign in1_94_10_ = ~(sub_844_2_n_151 ^ sub_844_2_n_11);
 assign sub_844_2_n_36 = ~(sub_844_2_n_117 | ~sub_844_2_n_142);
 assign sub_844_2_n_35 = ~(sub_844_2_n_121 | ~sub_844_2_n_122);
 assign in1_94_16_ = ~(sub_844_2_n_153 ^ sub_844_2_n_7);
 assign in1_94_8_ = (sub_844_2_n_146 ^ sub_844_2_n_4);
 assign in1_94_23_ = (sub_844_2_n_171 ^ sub_844_2_n_9);
 assign in1_94_9_ = (sub_844_2_n_150 ^ sub_844_2_n_108);
 assign in1_94_6_ = ~(sub_844_2_n_36 ^ sub_844_2_n_12);
 assign in1_94_22_ = ~(sub_844_2_n_169 ^ sub_844_2_n_3);
 assign in1_94_21_ = (sub_844_2_n_168 ^ sub_844_2_n_10);
 assign in1_94_2_ = (sub_844_2_n_135 ^ sub_844_2_n_103);
 assign in1_94_17_ = (sub_844_2_n_160 ^ sub_844_2_n_16);
 assign in1_94_11_ = (sub_844_2_n_157 ^ sub_844_2_n_98);
 assign sub_844_2_n_24 = ~(sub_844_2_n_112 | ~sub_844_2_n_97);
 assign in1_94_3_ = ~(sub_844_2_n_140 ^ sub_844_2_n_95);
 assign in1_94_13_ = (sub_844_2_n_158 ^ sub_844_2_n_17);
 assign in1_94_5_ = ~(sub_844_2_n_144 ^ sub_844_2_n_8);
 assign sub_844_2_n_20 = ~(sub_844_2_n_153 | ~sub_844_2_n_94);
 assign in1_94_12_ = (sub_844_2_n_152 ^ sub_844_2_n_14);
 assign in1_94_15_ = (sub_844_2_n_166 ^ sub_844_2_n_93);
 assign sub_844_2_n_17 = ~(sub_844_2_n_59 | ~sub_844_2_n_85);
 assign sub_844_2_n_16 = ~(sub_844_2_n_67 | ~sub_844_2_n_83);
 assign sub_844_2_n_15 = ~(sub_844_2_n_65 | ~sub_844_2_n_82);
 assign sub_844_2_n_14 = ~(sub_844_2_n_70 | ~sub_844_2_n_77);
 assign sub_844_2_n_13 = (sub_844_2_n_76 | sub_844_2_n_80);
 assign sub_844_2_n_12 = ~(sub_844_2_n_80 | ~sub_844_2_n_74);
 assign sub_844_2_n_11 = ~(sub_844_2_n_2 | ~sub_844_2_n_72);
 assign sub_844_2_n_10 = ~(sub_844_2_n_66 | ~sub_844_2_n_63);
 assign sub_844_2_n_9 = ~(sub_844_2_n_81 | ~sub_844_2_n_61);
 assign sub_844_2_n_8 = ~(sub_844_2_n_53 | ~sub_844_2_n_60);
 assign sub_844_2_n_7 = ~(sub_844_2_n_49 | ~sub_844_2_n_58);
 assign sub_844_2_n_6 = ~(sub_844_2_n_73 | ~sub_844_2_n_57);
 assign sub_844_2_n_5 = ~(sub_844_2_n_56 & ~sub_844_2_n_51);
 assign sub_844_2_n_4 = ~(sub_844_2_n_75 | ~sub_844_2_n_50);
 assign sub_844_2_n_3 = ~(sub_844_2_n_69 | ~sub_844_2_n_46);
 assign sub_844_2_n_2 = ~(in1_92_9_ | ~n_1551);
 assign sub_844_2_n_1 = ~(in1_92_2_ | ~n_1579);
 assign sub_844_2_n_0 = ~(in1_92_10_ | ~n_1555);
 assign sub_865_2_n_168 = ~(sub_865_2_n_63 & (sub_865_2_n_165 | sub_865_2_n_0));
 assign in1_97_21_ = ~(sub_865_2_n_163 ^ sub_865_2_n_97);
 assign in1_97_15_ = ~(sub_865_2_n_161 ^ sub_865_2_n_88);
 assign in1_97_24_ = (sub_865_2_n_156 ^ in1_95_23_);
 assign sub_865_2_n_163 = ~(sub_865_2_n_79 & (sub_865_2_n_157 | sub_865_2_n_6));
 assign sub_865_2_n_162 = ~(sub_865_2_n_54 & (sub_865_2_n_160 | sub_865_2_n_5));
 assign sub_865_2_n_161 = ~(sub_865_2_n_56 & (sub_865_2_n_159 | sub_865_2_n_59));
 assign sub_865_2_n_165 = ~(sub_865_2_n_109 | (sub_865_2_n_158 & sub_865_2_n_91));
 assign sub_865_2_n_158 = ~sub_865_2_n_157;
 assign sub_865_2_n_156 = ~(sub_865_2_n_134 | ((sub_865_2_n_146 & sub_865_2_n_122) | (sub_865_2_n_136
    & sub_865_2_n_122)));
 assign sub_865_2_n_155 = ~(sub_865_2_n_53 & (sub_865_2_n_150 | sub_865_2_n_2));
 assign sub_865_2_n_160 = ~(sub_865_2_n_43 | sub_865_2_n_110);
 assign sub_865_2_n_159 = ~(sub_865_2_n_111 | (sub_865_2_n_149 & sub_865_2_n_90));
 assign sub_865_2_n_157 = ~(sub_865_2_n_151 | sub_865_2_n_128);
 assign in1_97_16_ = ~(sub_865_2_n_150 ^ sub_865_2_n_10);
 assign sub_865_2_n_153 = ~(sub_865_2_n_58 & (sub_865_2_n_148 | sub_865_2_n_71));
 assign sub_865_2_n_152 = ~(sub_865_2_n_73 & (sub_865_2_n_44 | sub_865_2_n_75));
 assign sub_865_2_n_151 = ~(sub_865_2_n_150 | sub_865_2_n_117);
 assign sub_865_2_n_150 = ~(sub_865_2_n_146 | sub_865_2_n_136);
 assign sub_865_2_n_148 = ~sub_865_2_n_149;
 assign sub_865_2_n_149 = ~(sub_865_2_n_127 & (sub_865_2_n_144 | sub_865_2_n_39));
 assign sub_865_2_n_147 = ~(sub_865_2_n_51 & (sub_865_2_n_144 | sub_865_2_n_57));
 assign sub_865_2_n_146 = ~(sub_865_2_n_144 | sub_865_2_n_123);
 assign sub_865_2_n_145 = ~(sub_865_2_n_78 & (sub_865_2_n_143 | sub_865_2_n_1));
 assign sub_865_2_n_144 = ~(sub_865_2_n_126 | (sub_865_2_n_140 & sub_865_2_n_92));
 assign sub_865_2_n_143 = ~(sub_865_2_n_140 | sub_865_2_n_112);
 assign sub_865_2_n_142 = ~(sub_865_2_n_62 | (sub_865_2_n_137 & sub_865_2_n_64));
 assign in1_97_3_ = (sub_865_2_n_139 ^ sub_865_2_n_25);
 assign sub_865_2_n_140 = ~(sub_865_2_n_138 | sub_865_2_n_98);
 assign sub_865_2_n_139 = ~(sub_865_2_n_60 & (sub_865_2_n_133 | sub_865_2_n_74));
 assign sub_865_2_n_137 = ~sub_865_2_n_138;
 assign sub_865_2_n_138 = ~(sub_865_2_n_135 | sub_865_2_n_114);
 assign sub_865_2_n_136 = ~(sub_865_2_n_130 & (sub_865_2_n_127 | sub_865_2_n_121));
 assign sub_865_2_n_135 = ~(sub_865_2_n_133 | sub_865_2_n_22);
 assign sub_865_2_n_134 = ~(sub_865_2_n_129 & ~(sub_865_2_n_128 & sub_865_2_n_120));
 assign sub_865_2_n_133 = ~(sub_865_2_n_132 | sub_865_2_n_115);
 assign sub_865_2_n_132 = ~(sub_865_2_n_125 & ~(sub_865_2_n_70 & in1_95_0_));
 assign in1_97_1_ = (sub_865_2_n_116 ^ sub_865_2_n_70);
 assign sub_865_2_n_130 = ~(sub_865_2_n_105 | (sub_865_2_n_111 & sub_865_2_n_96));
 assign sub_865_2_n_129 = ~(sub_865_2_n_38 | sub_865_2_n_107);
 assign sub_865_2_n_128 = ~(sub_865_2_n_108 & ~(sub_865_2_n_110 & sub_865_2_n_100));
 assign sub_865_2_n_127 = ~(sub_865_2_n_124 | sub_865_2_n_113);
 assign sub_865_2_n_126 = ~(sub_865_2_n_106 & ~(sub_865_2_n_112 & sub_865_2_n_92));
 assign sub_865_2_n_125 = ~(sub_865_2_n_70 & ~n_1586);
 assign sub_865_2_n_124 = ~(sub_865_2_n_118 | sub_865_2_n_15);
 assign sub_865_2_n_123 = (sub_865_2_n_39 | sub_865_2_n_121);
 assign sub_865_2_n_122 = ~(sub_865_2_n_117 | sub_865_2_n_119);
 assign sub_865_2_n_120 = ~sub_865_2_n_119;
 assign sub_865_2_n_115 = (sub_865_2_n_49 & in1_95_0_);
 assign sub_865_2_n_116 = (sub_865_2_n_49 ^ in1_95_0_);
 assign sub_865_2_n_114 = ~(sub_865_2_n_83 & (sub_865_2_n_60 | sub_865_2_n_76));
 assign sub_865_2_n_113 = ~(sub_865_2_n_86 & (sub_865_2_n_73 | sub_865_2_n_8));
 assign sub_865_2_n_121 = ~(sub_865_2_n_90 & sub_865_2_n_96);
 assign sub_865_2_n_119 = ~(sub_865_2_n_91 & sub_865_2_n_103);
 assign sub_865_2_n_118 = ~(sub_865_2_n_82 | ~(sub_865_2_n_51 | sub_865_2_n_72));
 assign sub_865_2_n_117 = ~(sub_865_2_n_104 & sub_865_2_n_100);
 assign sub_865_2_n_108 = ~(sub_865_2_n_67 | ~(sub_865_2_n_54 | sub_865_2_n_80));
 assign sub_865_2_n_107 = ~(sub_865_2_n_68 & (sub_865_2_n_63 | sub_865_2_n_3));
 assign sub_865_2_n_106 = ~(sub_865_2_n_84 | ~(sub_865_2_n_78 | sub_865_2_n_52));
 assign sub_865_2_n_105 = ~(sub_865_2_n_66 & (sub_865_2_n_56 | sub_865_2_n_81));
 assign sub_865_2_n_112 = ~(sub_865_2_n_65 & (sub_865_2_n_61 | sub_865_2_n_77));
 assign sub_865_2_n_111 = ~(sub_865_2_n_87 & (sub_865_2_n_58 | sub_865_2_n_7));
 assign sub_865_2_n_110 = ~(sub_865_2_n_69 & (sub_865_2_n_53 | sub_865_2_n_4));
 assign sub_865_2_n_109 = ~(sub_865_2_n_85 & (sub_865_2_n_79 | sub_865_2_n_55));
 assign sub_865_2_n_98 = ~(sub_865_2_n_64 & ~sub_865_2_n_77);
 assign sub_865_2_n_104 = ~(sub_865_2_n_2 | sub_865_2_n_4);
 assign sub_865_2_n_103 = ~(sub_865_2_n_0 | sub_865_2_n_3);
 assign sub_865_2_n_102 = ~(sub_865_2_n_82 | sub_865_2_n_72);
 assign sub_865_2_n_97 = ~(sub_865_2_n_85 & ~sub_865_2_n_55);
 assign sub_865_2_n_101 = ~(sub_865_2_n_84 | sub_865_2_n_52);
 assign sub_865_2_n_100 = ~(sub_865_2_n_5 | sub_865_2_n_80);
 assign sub_865_2_n_99 = ~(sub_865_2_n_67 | sub_865_2_n_80);
 assign in1_97_0_ = ~(sub_865_2_n_70 & ~(sub_865_2_n_50 & n_1560));
 assign sub_865_2_n_96 = ~(sub_865_2_n_59 | sub_865_2_n_81);
 assign sub_865_2_n_95 = ~(sub_865_2_n_8 | ~sub_865_2_n_86);
 assign sub_865_2_n_94 = ~(sub_865_2_n_57 | sub_865_2_n_72);
 assign sub_865_2_n_93 = ~(sub_865_2_n_7 | ~sub_865_2_n_87);
 assign sub_865_2_n_92 = ~(sub_865_2_n_1 | sub_865_2_n_52);
 assign sub_865_2_n_88 = ~(sub_865_2_n_66 & ~sub_865_2_n_81);
 assign sub_865_2_n_91 = ~(sub_865_2_n_6 | sub_865_2_n_55);
 assign sub_865_2_n_90 = ~(sub_865_2_n_71 | sub_865_2_n_7);
 assign sub_865_2_n_87 = ~(in1_95_12_ & ~n_1581);
 assign sub_865_2_n_86 = ~(in1_95_10_ & ~n_1555);
 assign sub_865_2_n_85 = ~(in1_95_20_ & ~n_1593);
 assign sub_865_2_n_84 = ~(n_1527 | ~in1_95_6_);
 assign sub_865_2_n_83 = ~(in1_95_2_ & ~n_1579);
 assign sub_865_2_n_82 = ~(n_1589 | ~in1_95_8_);
 assign sub_865_2_n_81 = ~(in1_95_14_ | ~n_1495);
 assign sub_865_2_n_80 = ~(in1_95_18_ | ~n_1558);
 assign sub_865_2_n_79 = ~(in1_95_19_ & ~n_1565);
 assign sub_865_2_n_78 = ~(in1_95_5_ & ~n_1567);
 assign sub_865_2_n_77 = ~(in1_95_4_ | ~n_1569);
 assign sub_865_2_n_76 = ~(in1_95_2_ | ~n_1579);
 assign sub_865_2_n_75 = ~(in1_95_9_ | ~n_1551);
 assign sub_865_2_n_74 = ~(in1_95_1_ | ~n_1477);
 assign sub_865_2_n_73 = ~(in1_95_9_ & ~n_1551);
 assign sub_865_2_n_72 = ~(in1_95_8_ | ~n_1589);
 assign sub_865_2_n_71 = ~(in1_95_11_ | ~n_1595);
 assign sub_865_2_n_70 = ~(n_1543 & ~n_1560);
 assign sub_865_2_n_62 = ~sub_865_2_n_61;
 assign sub_865_2_n_69 = ~(in1_95_16_ & ~n_1562);
 assign sub_865_2_n_68 = ~(in1_95_22_ & ~n_1403);
 assign sub_865_2_n_67 = ~(n_1558 | ~in1_95_18_);
 assign sub_865_2_n_66 = ~(in1_95_14_ & ~n_1495);
 assign sub_865_2_n_65 = ~(in1_95_4_ & ~n_1569);
 assign sub_865_2_n_64 = ~(n_1535 & ~in1_95_3_);
 assign sub_865_2_n_63 = ~(in1_95_21_ & ~n_1591);
 assign sub_865_2_n_61 = ~(in1_95_3_ & ~n_1535);
 assign sub_865_2_n_60 = ~(in1_95_1_ & ~n_1477);
 assign sub_865_2_n_59 = ~(in1_95_13_ | ~n_1577);
 assign sub_865_2_n_58 = ~(in1_95_11_ & ~n_1595);
 assign sub_865_2_n_57 = ~(in1_95_7_ | ~n_1479);
 assign sub_865_2_n_56 = ~(in1_95_13_ & ~n_1577);
 assign sub_865_2_n_55 = ~(in1_95_20_ | ~n_1593);
 assign sub_865_2_n_54 = ~(in1_95_17_ & ~n_1472);
 assign sub_865_2_n_53 = ~(in1_95_15_ & ~n_1549);
 assign sub_865_2_n_52 = ~(in1_95_6_ | ~n_1527);
 assign sub_865_2_n_51 = ~(in1_95_7_ & ~n_1479);
 assign sub_865_2_n_50 = ~n_1543;
 assign sub_865_2_n_49 = ~n_1586;
 assign in1_97_18_ = ~(sub_865_2_n_160 ^ sub_865_2_n_11);
 assign in1_97_14_ = ~(sub_865_2_n_159 ^ sub_865_2_n_12);
 assign in1_97_10_ = ~(sub_865_2_n_44 ^ sub_865_2_n_21);
 assign in1_97_8_ = ~(sub_865_2_n_144 ^ sub_865_2_n_9);
 assign sub_865_2_n_44 = ~(sub_865_2_n_27 | ~sub_865_2_n_118);
 assign sub_865_2_n_43 = ~(sub_865_2_n_150 | ~sub_865_2_n_104);
 assign in1_97_6_ = ~(sub_865_2_n_143 ^ sub_865_2_n_23);
 assign in1_97_5_ = ~(sub_865_2_n_142 ^ sub_865_2_n_18);
 assign in1_97_2_ = ~(sub_865_2_n_133 ^ sub_865_2_n_14);
 assign sub_865_2_n_39 = ~(sub_865_2_n_94 & ~sub_865_2_n_15);
 assign sub_865_2_n_38 = (sub_865_2_n_103 & sub_865_2_n_109);
 assign in1_97_23_ = (sub_865_2_n_168 ^ sub_865_2_n_19);
 assign in1_97_9_ = (sub_865_2_n_147 ^ sub_865_2_n_102);
 assign in1_97_22_ = ~(sub_865_2_n_165 ^ sub_865_2_n_16);
 assign in1_97_7_ = (sub_865_2_n_145 ^ sub_865_2_n_101);
 assign in1_97_20_ = (sub_865_2_n_158 ^ sub_865_2_n_24);
 assign in1_97_19_ = (sub_865_2_n_162 ^ sub_865_2_n_99);
 assign in1_97_4_ = ~(sub_865_2_n_138 ^ sub_865_2_n_17);
 assign in1_97_17_ = (sub_865_2_n_155 ^ sub_865_2_n_20);
 assign in1_97_11_ = (sub_865_2_n_152 ^ sub_865_2_n_95);
 assign in1_97_12_ = (sub_865_2_n_149 ^ sub_865_2_n_13);
 assign sub_865_2_n_27 = ~(sub_865_2_n_144 | ~sub_865_2_n_94);
 assign in1_97_13_ = (sub_865_2_n_153 ^ sub_865_2_n_93);
 assign sub_865_2_n_25 = ~(sub_865_2_n_76 | ~sub_865_2_n_83);
 assign sub_865_2_n_24 = ~(sub_865_2_n_6 | ~sub_865_2_n_79);
 assign sub_865_2_n_23 = ~(sub_865_2_n_1 | ~sub_865_2_n_78);
 assign sub_865_2_n_22 = (sub_865_2_n_76 | sub_865_2_n_74);
 assign sub_865_2_n_21 = ~(sub_865_2_n_75 | ~sub_865_2_n_73);
 assign sub_865_2_n_20 = ~(sub_865_2_n_4 | ~sub_865_2_n_69);
 assign sub_865_2_n_19 = ~(sub_865_2_n_3 | ~sub_865_2_n_68);
 assign sub_865_2_n_18 = ~(sub_865_2_n_77 | ~sub_865_2_n_65);
 assign sub_865_2_n_17 = ~(sub_865_2_n_62 | ~sub_865_2_n_64);
 assign sub_865_2_n_16 = ~(sub_865_2_n_0 | ~sub_865_2_n_63);
 assign sub_865_2_n_15 = (sub_865_2_n_8 | sub_865_2_n_75);
 assign sub_865_2_n_14 = ~(sub_865_2_n_74 | ~sub_865_2_n_60);
 assign sub_865_2_n_13 = ~(sub_865_2_n_71 | ~sub_865_2_n_58);
 assign sub_865_2_n_12 = ~(sub_865_2_n_59 | ~sub_865_2_n_56);
 assign sub_865_2_n_11 = ~(sub_865_2_n_5 | ~sub_865_2_n_54);
 assign sub_865_2_n_10 = ~(sub_865_2_n_2 | ~sub_865_2_n_53);
 assign sub_865_2_n_9 = ~(sub_865_2_n_57 | ~sub_865_2_n_51);
 assign sub_865_2_n_8 = ~(in1_95_10_ | ~n_1555);
 assign sub_865_2_n_7 = ~(in1_95_12_ | ~n_1581);
 assign sub_865_2_n_6 = ~(in1_95_19_ | ~n_1565);
 assign sub_865_2_n_5 = ~(in1_95_17_ | ~n_1472);
 assign sub_865_2_n_4 = ~(in1_95_16_ | ~n_1562);
 assign sub_865_2_n_3 = ~(in1_95_22_ | ~n_1403);
 assign sub_865_2_n_2 = ~(in1_95_15_ | ~n_1549);
 assign sub_865_2_n_1 = ~(in1_95_5_ | ~n_1567);
 assign sub_865_2_n_0 = ~(in1_95_21_ | ~n_1591);
 assign sub_886_2_n_178 = ~(sub_886_2_n_44 | (sub_886_2_n_177 & sub_886_2_n_71));
 assign sub_886_2_n_177 = ~(sub_886_2_n_123 & (sub_886_2_n_172 | sub_886_2_n_98));
 assign sub_886_2_n_176 = ~(sub_886_2_n_173 | sub_886_2_n_43);
 assign sub_886_2_n_175 = ~(sub_886_2_n_57 | (sub_886_2_n_171 & sub_886_2_n_3));
 assign sub_886_2_n_174 = ~(sub_886_2_n_81 & (sub_886_2_n_169 | sub_886_2_n_66));
 assign sub_886_2_n_173 = ~(sub_886_2_n_172 | sub_886_2_n_79);
 assign sub_886_2_n_172 = ~(sub_886_2_n_138 | ~(sub_886_2_n_162 | sub_886_2_n_27));
 assign sub_886_2_n_171 = ~(sub_886_2_n_122 & (sub_886_2_n_162 | sub_886_2_n_94));
 assign sub_886_2_n_170 = ~(sub_886_2_n_164 | sub_886_2_n_59);
 assign sub_886_2_n_169 = ~(sub_886_2_n_125 | (sub_886_2_n_160 & sub_886_2_n_110));
 assign sub_886_2_n_168 = ~(sub_886_2_n_78 & (sub_886_2_n_161 | sub_886_2_n_72));
 assign sub_886_2_n_167 = ~(sub_886_2_n_73 & (sub_886_2_n_33 | sub_886_2_n_47));
 assign in1_100_16_ = ~(sub_886_2_n_162 ^ sub_886_2_n_104);
 assign in1_100_12_ = ~(sub_886_2_n_160 ^ sub_886_2_n_88);
 assign sub_886_2_n_164 = ~(sub_886_2_n_162 | sub_886_2_n_46);
 assign sub_886_2_n_163 = ~(sub_886_2_n_150 | (sub_886_2_n_156 & sub_886_2_n_133));
 assign sub_886_2_n_162 = ~(sub_886_2_n_156 | sub_886_2_n_146);
 assign sub_886_2_n_161 = ~sub_886_2_n_160;
 assign sub_886_2_n_160 = ~(sub_886_2_n_141 & (sub_886_2_n_155 | sub_886_2_n_21));
 assign sub_886_2_n_159 = ~(sub_886_2_n_48 & (sub_886_2_n_155 | sub_886_2_n_76));
 assign in1_100_8_ = ~(sub_886_2_n_155 ^ sub_886_2_n_6);
 assign sub_886_2_n_157 = ~(sub_886_2_n_75 | (sub_886_2_n_153 & sub_886_2_n_0));
 assign sub_886_2_n_156 = ~(sub_886_2_n_155 | sub_886_2_n_135);
 assign sub_886_2_n_155 = ~(sub_886_2_n_154 | sub_886_2_n_140);
 assign sub_886_2_n_154 = ~(sub_886_2_n_151 | sub_886_2_n_116);
 assign sub_886_2_n_153 = ~(sub_886_2_n_151 & sub_886_2_n_126);
 assign sub_886_2_n_152 = ~(sub_886_2_n_50 | (sub_886_2_n_148 & sub_886_2_n_53));
 assign sub_886_2_n_151 = ~(sub_886_2_n_148 & sub_886_2_n_106);
 assign sub_886_2_n_150 = ~(sub_886_2_n_145 & ~(sub_886_2_n_146 & sub_886_2_n_133));
 assign sub_886_2_n_149 = ~(sub_886_2_n_40 & (sub_886_2_n_144 | sub_886_2_n_45));
 assign sub_886_2_n_148 = ~(sub_886_2_n_147 & sub_886_2_n_119);
 assign sub_886_2_n_147 = ~(sub_886_2_n_143 & sub_886_2_n_91);
 assign sub_886_2_n_146 = ~(sub_886_2_n_139 & (sub_886_2_n_141 | sub_886_2_n_30));
 assign sub_886_2_n_145 = ~(sub_886_2_n_137 | (sub_886_2_n_138 & sub_886_2_n_131));
 assign sub_886_2_n_144 = ~sub_886_2_n_143;
 assign sub_886_2_n_143 = ((sub_886_2_n_39 & in1_98_0_) | ((in1_98_0_ & sub_886_2_n_38) | (sub_886_2_n_38
    & sub_886_2_n_39)));
 assign in1_100_1_ = (in1_98_0_ ^ (sub_886_2_n_38 ^ sub_886_2_n_39));
 assign sub_886_2_n_141 = ~(sub_886_2_n_134 | sub_886_2_n_120);
 assign sub_886_2_n_140 = ~(sub_886_2_n_128 & (sub_886_2_n_126 | sub_886_2_n_116));
 assign sub_886_2_n_139 = ~(sub_886_2_n_136 | sub_886_2_n_129);
 assign sub_886_2_n_138 = ~(sub_886_2_n_127 & (sub_886_2_n_122 | sub_886_2_n_5));
 assign sub_886_2_n_137 = ~(sub_886_2_n_132 & sub_886_2_n_118);
 assign sub_886_2_n_136 = ~(sub_886_2_n_124 | sub_886_2_n_114);
 assign sub_886_2_n_135 = (sub_886_2_n_21 | sub_886_2_n_30);
 assign sub_886_2_n_134 = ~(sub_886_2_n_121 | sub_886_2_n_7);
 assign sub_886_2_n_133 = ~(sub_886_2_n_27 | sub_886_2_n_130);
 assign sub_886_2_n_132 = ~(sub_886_2_n_113 & ~sub_886_2_n_123);
 assign sub_886_2_n_131 = ~sub_886_2_n_130;
 assign sub_886_2_n_129 = ~(sub_886_2_n_63 & (sub_886_2_n_81 | sub_886_2_n_51));
 assign sub_886_2_n_128 = ~(sub_886_2_n_65 | ~(sub_886_2_n_74 | sub_886_2_n_77));
 assign sub_886_2_n_127 = ~(sub_886_2_n_86 | ~(sub_886_2_n_56 | sub_886_2_n_41));
 assign sub_886_2_n_130 = ~(sub_886_2_n_113 & ~sub_886_2_n_98);
 assign sub_886_2_n_125 = ~sub_886_2_n_124;
 assign sub_886_2_n_120 = ~(sub_886_2_n_85 & (sub_886_2_n_73 | sub_886_2_n_54));
 assign sub_886_2_n_119 = ~(sub_886_2_n_87 | ~(sub_886_2_n_40 | sub_886_2_n_55));
 assign sub_886_2_n_118 = ~(sub_886_2_n_90 | sub_886_2_n_62);
 assign sub_886_2_n_126 = ~(sub_886_2_n_107 | sub_886_2_n_61);
 assign sub_886_2_n_124 = ~(sub_886_2_n_84 | ~(sub_886_2_n_78 | sub_886_2_n_60));
 assign sub_886_2_n_123 = ~(sub_886_2_n_105 | sub_886_2_n_64);
 assign sub_886_2_n_122 = ~(sub_886_2_n_82 | ~(sub_886_2_n_58 | sub_886_2_n_68));
 assign sub_886_2_n_121 = ~(sub_886_2_n_83 | ~(sub_886_2_n_48 | sub_886_2_n_69));
 assign sub_886_2_n_107 = ~(sub_886_2_n_49 | sub_886_2_n_2);
 assign sub_886_2_n_106 = ~(sub_886_2_n_52 | sub_886_2_n_2);
 assign sub_886_2_n_105 = ~(sub_886_2_n_42 | sub_886_2_n_67);
 assign sub_886_2_n_117 = ~(sub_886_2_n_44 | sub_886_2_n_70);
 assign sub_886_2_n_116 = ~(sub_886_2_n_0 & ~sub_886_2_n_77);
 assign sub_886_2_n_115 = ~(sub_886_2_n_83 | sub_886_2_n_69);
 assign sub_886_2_n_114 = (sub_886_2_n_66 | sub_886_2_n_51);
 assign sub_886_2_n_113 = ~(sub_886_2_n_70 | sub_886_2_n_80);
 assign sub_886_2_n_112 = ~(sub_886_2_n_62 | sub_886_2_n_80);
 assign sub_886_2_n_111 = ~(sub_886_2_n_64 | sub_886_2_n_67);
 assign sub_886_2_n_110 = ~(sub_886_2_n_72 | sub_886_2_n_60);
 assign sub_886_2_n_109 = ~(sub_886_2_n_43 | sub_886_2_n_79);
 assign sub_886_2_n_108 = ~(sub_886_2_n_86 | sub_886_2_n_41);
 assign sub_886_2_n_104 = ~(sub_886_2_n_59 | sub_886_2_n_46);
 assign sub_886_2_n_94 = ~sub_886_2_n_93;
 assign sub_886_2_n_91 = ~(sub_886_2_n_45 | sub_886_2_n_55);
 assign sub_886_2_n_90 = ~(sub_886_2_n_80 | ~sub_886_2_n_44);
 assign in1_100_0_ = ~(sub_886_2_n_39 & ~(sub_886_2_n_37 & n_1564));
 assign sub_886_2_n_103 = ~(sub_886_2_n_82 | sub_886_2_n_68);
 assign sub_886_2_n_102 = ~(sub_886_2_n_54 | ~sub_886_2_n_85);
 assign sub_886_2_n_101 = ~(sub_886_2_n_76 | sub_886_2_n_69);
 assign sub_886_2_n_100 = ~(sub_886_2_n_87 | sub_886_2_n_55);
 assign sub_886_2_n_99 = ~(sub_886_2_n_51 | ~sub_886_2_n_63);
 assign sub_886_2_n_98 = (sub_886_2_n_79 | sub_886_2_n_67);
 assign sub_886_2_n_97 = ~(sub_886_2_n_65 | sub_886_2_n_77);
 assign sub_886_2_n_96 = ~(sub_886_2_n_84 | sub_886_2_n_60);
 assign sub_886_2_n_95 = ~(sub_886_2_n_61 | sub_886_2_n_2);
 assign sub_886_2_n_93 = ~(sub_886_2_n_46 | sub_886_2_n_68);
 assign sub_886_2_n_88 = ~(sub_886_2_n_78 & ~sub_886_2_n_72);
 assign sub_886_2_n_92 = ~(sub_886_2_n_50 | sub_886_2_n_52);
 assign sub_886_2_n_75 = ~sub_886_2_n_74;
 assign sub_886_2_n_71 = ~sub_886_2_n_70;
 assign sub_886_2_n_87 = ~(n_1579 | ~in1_98_2_);
 assign sub_886_2_n_86 = ~(n_1558 | ~in1_98_18_);
 assign sub_886_2_n_85 = ~(in1_98_10_ & ~n_1555);
 assign sub_886_2_n_84 = ~(n_1581 | ~in1_98_12_);
 assign sub_886_2_n_83 = ~(n_1589 | ~in1_98_8_);
 assign sub_886_2_n_82 = ~(n_1562 | ~in1_98_16_);
 assign sub_886_2_n_81 = ~(in1_98_13_ & ~n_1577);
 assign sub_886_2_n_80 = ~(in1_98_22_ | sub_886_2_n_36);
 assign sub_886_2_n_79 = ~(in1_98_19_ | ~n_1565);
 assign sub_886_2_n_78 = ~(in1_98_11_ & ~n_1595);
 assign sub_886_2_n_77 = ~(in1_98_6_ | ~n_1527);
 assign sub_886_2_n_76 = ~(in1_98_7_ | ~n_1479);
 assign sub_886_2_n_74 = ~(in1_98_5_ & ~n_1567);
 assign sub_886_2_n_73 = ~(in1_98_9_ & ~n_1551);
 assign sub_886_2_n_72 = ~(in1_98_11_ | ~n_1595);
 assign sub_886_2_n_70 = ~(in1_98_21_ | ~n_1591);
 assign sub_886_2_n_69 = ~(in1_98_8_ | ~n_1589);
 assign sub_886_2_n_68 = ~(in1_98_16_ | ~n_1562);
 assign sub_886_2_n_67 = ~(in1_98_20_ | ~n_1593);
 assign sub_886_2_n_66 = ~(in1_98_13_ | ~n_1577);
 assign sub_886_2_n_59 = ~sub_886_2_n_58;
 assign sub_886_2_n_57 = ~sub_886_2_n_56;
 assign sub_886_2_n_53 = ~sub_886_2_n_52;
 assign sub_886_2_n_50 = ~sub_886_2_n_49;
 assign sub_886_2_n_43 = ~sub_886_2_n_42;
 assign sub_886_2_n_65 = ~(n_1527 | ~in1_98_6_);
 assign sub_886_2_n_64 = ~(n_1593 | ~in1_98_20_);
 assign sub_886_2_n_63 = ~(in1_98_14_ & ~n_1495);
 assign sub_886_2_n_62 = (sub_886_2_n_36 & in1_98_22_);
 assign sub_886_2_n_61 = ~(n_1569 | ~in1_98_4_);
 assign sub_886_2_n_60 = ~(in1_98_12_ | ~n_1581);
 assign sub_886_2_n_58 = ~(in1_98_15_ & ~n_1549);
 assign sub_886_2_n_56 = ~(in1_98_17_ & ~n_1472);
 assign sub_886_2_n_55 = ~(in1_98_2_ | ~n_1579);
 assign sub_886_2_n_54 = ~(in1_98_10_ | ~n_1555);
 assign sub_886_2_n_52 = ~(in1_98_3_ | ~n_1535);
 assign sub_886_2_n_51 = ~(in1_98_14_ | ~n_1495);
 assign sub_886_2_n_49 = ~(in1_98_3_ & ~n_1535);
 assign sub_886_2_n_48 = ~(in1_98_7_ & ~n_1479);
 assign sub_886_2_n_47 = ~(in1_98_9_ | ~n_1551);
 assign sub_886_2_n_46 = ~(in1_98_15_ | ~n_1549);
 assign sub_886_2_n_45 = ~(in1_98_1_ | ~n_1477);
 assign sub_886_2_n_44 = ~(n_1591 | ~in1_98_21_);
 assign sub_886_2_n_42 = ~(in1_98_19_ & ~n_1565);
 assign sub_886_2_n_41 = ~(in1_98_18_ | ~n_1558);
 assign sub_886_2_n_40 = ~(in1_98_1_ & ~n_1477);
 assign sub_886_2_n_39 = ~(n_1543 & ~n_1564);
 assign sub_886_2_n_38 = ~n_1586;
 assign sub_886_2_n_37 = ~n_1543;
 assign sub_886_2_n_36 = ~n_1403;
 assign in1_100_18_ = (sub_886_2_n_171 ^ sub_886_2_n_9);
 assign in1_100_6_ = (sub_886_2_n_153 ^ sub_886_2_n_10);
 assign sub_886_2_n_33 = ~(sub_886_2_n_20 | ~sub_886_2_n_121);
 assign in1_100_22_ = (sub_886_2_n_177 ^ sub_886_2_n_117);
 assign in1_100_9_ = (sub_886_2_n_159 ^ sub_886_2_n_115);
 assign sub_886_2_n_30 = ~(sub_886_2_n_110 & ~sub_886_2_n_114);
 assign in1_100_23_ = ~(sub_886_2_n_178 ^ sub_886_2_n_112);
 assign in1_100_21_ = ~(sub_886_2_n_176 ^ sub_886_2_n_111);
 assign sub_886_2_n_27 = ~(sub_886_2_n_93 & ~sub_886_2_n_5);
 assign in1_100_20_ = ~(sub_886_2_n_172 ^ sub_886_2_n_109);
 assign in1_100_2_ = (sub_886_2_n_143 ^ sub_886_2_n_4);
 assign in1_100_19_ = ~(sub_886_2_n_175 ^ sub_886_2_n_108);
 assign in1_100_17_ = ~(sub_886_2_n_170 ^ sub_886_2_n_103);
 assign in1_100_11_ = (sub_886_2_n_167 ^ sub_886_2_n_102);
 assign sub_886_2_n_21 = ~(sub_886_2_n_101 & ~sub_886_2_n_7);
 assign sub_886_2_n_20 = ~(sub_886_2_n_155 | ~sub_886_2_n_101);
 assign in1_100_3_ = (sub_886_2_n_149 ^ sub_886_2_n_100);
 assign in1_100_15_ = (sub_886_2_n_174 ^ sub_886_2_n_99);
 assign in1_100_7_ = ~(sub_886_2_n_157 ^ sub_886_2_n_97);
 assign in1_100_14_ = ~(sub_886_2_n_169 ^ sub_886_2_n_11);
 assign in1_100_13_ = (sub_886_2_n_168 ^ sub_886_2_n_96);
 assign in1_100_5_ = ~(sub_886_2_n_152 ^ sub_886_2_n_95);
 assign in1_100_10_ = ~(sub_886_2_n_33 ^ sub_886_2_n_8);
 assign in1_100_4_ = (sub_886_2_n_148 ^ sub_886_2_n_92);
 assign sub_886_2_n_11 = ~(sub_886_2_n_66 | ~sub_886_2_n_81);
 assign sub_886_2_n_10 = ~(sub_886_2_n_75 | ~sub_886_2_n_0);
 assign sub_886_2_n_9 = ~(sub_886_2_n_57 | ~sub_886_2_n_3);
 assign sub_886_2_n_8 = ~(sub_886_2_n_47 | ~sub_886_2_n_73);
 assign sub_886_2_n_7 = (sub_886_2_n_54 | sub_886_2_n_47);
 assign sub_886_2_n_6 = ~(sub_886_2_n_76 | ~sub_886_2_n_48);
 assign sub_886_2_n_5 = ~(sub_886_2_n_3 & ~sub_886_2_n_41);
 assign sub_886_2_n_4 = ~(sub_886_2_n_45 | ~sub_886_2_n_40);
 assign sub_886_2_n_3 = ~(n_1472 & ~in1_98_17_);
 assign sub_886_2_n_2 = ~(in1_98_4_ | ~n_1569);
 assign in1_100_24_ = (sub_886_2_n_163 ^ in1_98_23_);
 assign sub_886_2_n_0 = ~(n_1567 & ~in1_98_5_);
 assign sub_907_2_n_169 = ~(sub_907_2_n_46 & (sub_907_2_n_167 | sub_907_2_n_44));
 assign in1_103_21_ = ~(sub_907_2_n_165 ^ sub_907_2_n_17);
 assign sub_907_2_n_167 = ~sub_907_2_n_166;
 assign sub_907_2_n_166 = ~(sub_907_2_n_109 & (sub_907_2_n_161 | sub_907_2_n_89));
 assign sub_907_2_n_165 = ~(sub_907_2_n_69 & (sub_907_2_n_161 | sub_907_2_n_68));
 assign sub_907_2_n_164 = ~(sub_907_2_n_74 & (sub_907_2_n_160 | sub_907_2_n_48));
 assign sub_907_2_n_163 = ~(sub_907_2_n_42 & (sub_907_2_n_154 | sub_907_2_n_41));
 assign in1_103_24_ = ~(sub_907_2_n_155 ^ in1_101_23_);
 assign sub_907_2_n_161 = ~(sub_907_2_n_156 | sub_907_2_n_126);
 assign sub_907_2_n_160 = ~(sub_907_2_n_20 | sub_907_2_n_110);
 assign sub_907_2_n_159 = ~(sub_907_2_n_72 & (sub_907_2_n_34 | sub_907_2_n_3));
 assign in1_103_16_ = (sub_907_2_n_34 ^ sub_907_2_n_83);
 assign in1_103_11_ = ~(sub_907_2_n_150 ^ sub_907_2_n_93);
 assign sub_907_2_n_156 = ~(sub_907_2_n_34 | sub_907_2_n_113);
 assign sub_907_2_n_155 = ~(sub_907_2_n_134 & (sub_907_2_n_148 | sub_907_2_n_118));
 assign sub_907_2_n_154 = ~(sub_907_2_n_151 | sub_907_2_n_114);
 assign sub_907_2_n_153 = ~(sub_907_2_n_73 & (sub_907_2_n_147 | sub_907_2_n_49));
 assign in1_103_12_ = (sub_907_2_n_147 ^ sub_907_2_n_82);
 assign sub_907_2_n_151 = ~(sub_907_2_n_147 | sub_907_2_n_99);
 assign sub_907_2_n_150 = ~(sub_907_2_n_65 & (sub_907_2_n_33 | sub_907_2_n_43));
 assign in1_103_10_ = (sub_907_2_n_33 ^ sub_907_2_n_86);
 assign sub_907_2_n_148 = ~(sub_907_2_n_23 & sub_907_2_n_29);
 assign sub_907_2_n_147 = ~(sub_907_2_n_23 | sub_907_2_n_124);
 assign in1_103_7_ = (sub_907_2_n_143 ^ sub_907_2_n_85);
 assign sub_907_2_n_145 = ~(sub_907_2_n_40 & (sub_907_2_n_141 | sub_907_2_n_50));
 assign in1_103_8_ = ~(sub_907_2_n_141 ^ sub_907_2_n_4);
 assign sub_907_2_n_143 = ~(sub_907_2_n_67 & (sub_907_2_n_139 | sub_907_2_n_61));
 assign sub_907_2_n_142 = ~(sub_907_2_n_140 & sub_907_2_n_88);
 assign sub_907_2_n_141 = ~sub_907_2_n_140;
 assign sub_907_2_n_140 = ~(sub_907_2_n_138 & sub_907_2_n_125);
 assign sub_907_2_n_139 = ~(sub_907_2_n_135 | sub_907_2_n_108);
 assign sub_907_2_n_138 = ~(sub_907_2_n_135 & sub_907_2_n_101);
 assign sub_907_2_n_137 = ~(sub_907_2_n_70 | (sub_907_2_n_131 & sub_907_2_n_63));
 assign in1_103_3_ = (sub_907_2_n_132 ^ sub_907_2_n_84);
 assign sub_907_2_n_135 = ~(sub_907_2_n_130 | sub_907_2_n_95);
 assign sub_907_2_n_134 = ~(sub_907_2_n_133 | sub_907_2_n_127);
 assign sub_907_2_n_133 = ~(sub_907_2_n_128 | sub_907_2_n_118);
 assign sub_907_2_n_132 = ~(sub_907_2_n_47 & (sub_907_2_n_121 | sub_907_2_n_66));
 assign sub_907_2_n_131 = ~sub_907_2_n_130;
 assign sub_907_2_n_130 = ~(sub_907_2_n_129 | sub_907_2_n_105);
 assign sub_907_2_n_129 = ~(sub_907_2_n_121 | sub_907_2_n_15);
 assign sub_907_2_n_128 = ~(sub_907_2_n_123 | (sub_907_2_n_124 & sub_907_2_n_29));
 assign sub_907_2_n_127 = ~(sub_907_2_n_122 & ~(sub_907_2_n_126 & sub_907_2_n_116));
 assign sub_907_2_n_126 = ~(sub_907_2_n_106 & ~(sub_907_2_n_110 & sub_907_2_n_98));
 assign sub_907_2_n_125 = ~(sub_907_2_n_107 | (sub_907_2_n_108 & sub_907_2_n_101));
 assign sub_907_2_n_124 = ~(sub_907_2_n_120 & sub_907_2_n_111);
 assign sub_907_2_n_123 = ~(sub_907_2_n_112 & ~(sub_907_2_n_114 & sub_907_2_n_102));
 assign sub_907_2_n_122 = ~(sub_907_2_n_119 | sub_907_2_n_104);
 assign sub_907_2_n_121 = ~(sub_907_2_n_117 | sub_907_2_n_56);
 assign sub_907_2_n_120 = ~(sub_907_2_n_115 & sub_907_2_n_92);
 assign sub_907_2_n_119 = ~(sub_907_2_n_109 | sub_907_2_n_100);
 assign sub_907_2_n_118 = ~(sub_907_2_n_116 & ~sub_907_2_n_113);
 assign sub_907_2_n_117 = ~(sub_907_2_n_57 | ~sub_907_2_n_39);
 assign sub_907_2_n_112 = ~(sub_907_2_n_54 | ~(sub_907_2_n_42 | sub_907_2_n_64));
 assign sub_907_2_n_111 = ~(sub_907_2_n_80 | ~(sub_907_2_n_65 | sub_907_2_n_51));
 assign sub_907_2_n_116 = ~(sub_907_2_n_89 | sub_907_2_n_100);
 assign sub_907_2_n_115 = ~(sub_907_2_n_58 & (sub_907_2_n_40 | sub_907_2_n_0));
 assign sub_907_2_n_114 = ~(sub_907_2_n_55 & (sub_907_2_n_73 | sub_907_2_n_45));
 assign sub_907_2_n_113 = ~(sub_907_2_n_90 & sub_907_2_n_98);
 assign sub_907_2_n_107 = ~(sub_907_2_n_78 & (sub_907_2_n_67 | sub_907_2_n_62));
 assign sub_907_2_n_106 = ~(sub_907_2_n_77 | ~(sub_907_2_n_74 | sub_907_2_n_52));
 assign sub_907_2_n_105 = ~(sub_907_2_n_76 & (sub_907_2_n_47 | sub_907_2_n_75));
 assign sub_907_2_n_104 = ~(sub_907_2_n_53 & (sub_907_2_n_46 | sub_907_2_n_71));
 assign sub_907_2_n_110 = ~(sub_907_2_n_79 & (sub_907_2_n_72 | sub_907_2_n_1));
 assign sub_907_2_n_109 = ~(sub_907_2_n_81 | ~(sub_907_2_n_69 | sub_907_2_n_60));
 assign sub_907_2_n_108 = ~(sub_907_2_n_96 & sub_907_2_n_59);
 assign sub_907_2_n_96 = ~(sub_907_2_n_70 & sub_907_2_n_2);
 assign sub_907_2_n_95 = ~(sub_907_2_n_63 & sub_907_2_n_2);
 assign sub_907_2_n_94 = ~(sub_907_2_n_56 | sub_907_2_n_57);
 assign sub_907_2_n_103 = ~(sub_907_2_n_71 | ~sub_907_2_n_53);
 assign sub_907_2_n_102 = ~(sub_907_2_n_41 | sub_907_2_n_64);
 assign sub_907_2_n_101 = ~(sub_907_2_n_61 | sub_907_2_n_62);
 assign sub_907_2_n_100 = (sub_907_2_n_44 | sub_907_2_n_71);
 assign sub_907_2_n_93 = (sub_907_2_n_80 | sub_907_2_n_51);
 assign sub_907_2_n_99 = (sub_907_2_n_49 | sub_907_2_n_45);
 assign sub_907_2_n_98 = ~(sub_907_2_n_48 | sub_907_2_n_52);
 assign sub_907_2_n_97 = ~(sub_907_2_n_77 | sub_907_2_n_52);
 assign sub_907_2_n_88 = ~(sub_907_2_n_50 | sub_907_2_n_0);
 assign in1_103_0_ = ~(sub_907_2_n_39 & ~(sub_907_2_n_38 & n_1548));
 assign sub_907_2_n_86 = ~(sub_907_2_n_65 & ~sub_907_2_n_43);
 assign sub_907_2_n_92 = ~(sub_907_2_n_43 | sub_907_2_n_51);
 assign sub_907_2_n_85 = ~(sub_907_2_n_62 | ~sub_907_2_n_78);
 assign sub_907_2_n_84 = ~(sub_907_2_n_75 | ~sub_907_2_n_76);
 assign sub_907_2_n_91 = ~(sub_907_2_n_54 | sub_907_2_n_64);
 assign sub_907_2_n_83 = ~(sub_907_2_n_72 & ~sub_907_2_n_3);
 assign sub_907_2_n_82 = ~(sub_907_2_n_73 & ~sub_907_2_n_49);
 assign sub_907_2_n_90 = ~(sub_907_2_n_3 | sub_907_2_n_1);
 assign sub_907_2_n_89 = (sub_907_2_n_68 | sub_907_2_n_60);
 assign sub_907_2_n_81 = ~(n_1593 | ~in1_101_20_);
 assign sub_907_2_n_80 = ~(n_1555 | ~in1_101_10_);
 assign sub_907_2_n_79 = ~(in1_101_16_ & ~n_1562);
 assign sub_907_2_n_78 = ~(in1_101_6_ & ~n_1527);
 assign sub_907_2_n_77 = ~(n_1558 | ~in1_101_18_);
 assign sub_907_2_n_76 = ~(in1_101_2_ & ~n_1579);
 assign sub_907_2_n_75 = ~(in1_101_2_ | ~n_1579);
 assign sub_907_2_n_74 = ~(in1_101_17_ & ~n_1472);
 assign sub_907_2_n_73 = ~(in1_101_11_ & ~n_1595);
 assign sub_907_2_n_72 = ~(in1_101_15_ & ~n_1549);
 assign sub_907_2_n_71 = ~(in1_101_22_ | ~n_1403);
 assign sub_907_2_n_70 = ~(n_1535 | ~in1_101_3_);
 assign sub_907_2_n_69 = ~(in1_101_19_ & ~n_1565);
 assign sub_907_2_n_68 = ~(in1_101_19_ | ~n_1565);
 assign sub_907_2_n_67 = ~(in1_101_5_ & ~n_1567);
 assign sub_907_2_n_66 = ~(in1_101_1_ | ~n_1477);
 assign sub_907_2_n_65 = ~(in1_101_9_ & ~n_1551);
 assign sub_907_2_n_64 = ~(in1_101_14_ | ~n_1495);
 assign sub_907_2_n_63 = ~(n_1535 & ~in1_101_3_);
 assign sub_907_2_n_62 = ~(in1_101_6_ | ~n_1527);
 assign sub_907_2_n_61 = ~(in1_101_5_ | ~n_1567);
 assign sub_907_2_n_60 = ~(in1_101_20_ | ~n_1593);
 assign sub_907_2_n_59 = ~(in1_101_4_ & ~n_1569);
 assign sub_907_2_n_58 = ~(in1_101_8_ & ~n_1589);
 assign sub_907_2_n_57 = ~(in1_101_0_ | ~n_1586);
 assign sub_907_2_n_56 = ~(n_1586 | ~in1_101_0_);
 assign sub_907_2_n_55 = ~(in1_101_12_ & ~n_1581);
 assign sub_907_2_n_54 = ~(n_1495 | ~in1_101_14_);
 assign sub_907_2_n_53 = ~(in1_101_22_ & ~n_1403);
 assign sub_907_2_n_52 = ~(in1_101_18_ | ~n_1558);
 assign sub_907_2_n_51 = ~(in1_101_10_ | ~n_1555);
 assign sub_907_2_n_50 = ~(in1_101_7_ | ~n_1479);
 assign sub_907_2_n_49 = ~(in1_101_11_ | ~n_1595);
 assign sub_907_2_n_48 = ~(in1_101_17_ | ~n_1472);
 assign sub_907_2_n_47 = ~(in1_101_1_ & ~n_1477);
 assign sub_907_2_n_46 = ~(in1_101_21_ & ~n_1591);
 assign sub_907_2_n_45 = ~(in1_101_12_ | ~n_1581);
 assign sub_907_2_n_44 = ~(in1_101_21_ | ~n_1591);
 assign sub_907_2_n_43 = ~(in1_101_9_ | ~n_1551);
 assign sub_907_2_n_42 = ~(in1_101_13_ & ~n_1577);
 assign sub_907_2_n_41 = ~(in1_101_13_ | ~n_1577);
 assign sub_907_2_n_40 = ~(in1_101_7_ & ~n_1479);
 assign sub_907_2_n_39 = ~(n_1543 & ~n_1548);
 assign sub_907_2_n_38 = ~n_1543;
 assign in1_103_20_ = ~(sub_907_2_n_161 ^ sub_907_2_n_13);
 assign in1_103_18_ = ~(sub_907_2_n_160 ^ sub_907_2_n_14);
 assign in1_103_14_ = ~(sub_907_2_n_154 ^ sub_907_2_n_5);
 assign sub_907_2_n_34 = (sub_907_2_n_148 & sub_907_2_n_128);
 assign sub_907_2_n_33 = ~(sub_907_2_n_115 | ~sub_907_2_n_142);
 assign in1_103_2_ = ~(sub_907_2_n_121 ^ sub_907_2_n_7);
 assign in1_103_1_ = (sub_907_2_n_94 ^ sub_907_2_n_39);
 assign in1_103_23_ = (sub_907_2_n_169 ^ sub_907_2_n_103);
 assign sub_907_2_n_29 = ~(sub_907_2_n_99 | ~sub_907_2_n_102);
 assign in1_103_5_ = ~(sub_907_2_n_137 ^ sub_907_2_n_10);
 assign in1_103_22_ = (sub_907_2_n_166 ^ sub_907_2_n_6);
 assign in1_103_6_ = ~(sub_907_2_n_139 ^ sub_907_2_n_12);
 assign in1_103_19_ = (sub_907_2_n_164 ^ sub_907_2_n_97);
 assign in1_103_4_ = ~(sub_907_2_n_130 ^ sub_907_2_n_11);
 assign sub_907_2_n_23 = ~(sub_907_2_n_142 | ~sub_907_2_n_92);
 assign in1_103_15_ = (sub_907_2_n_163 ^ sub_907_2_n_91);
 assign in1_103_13_ = (sub_907_2_n_153 ^ sub_907_2_n_8);
 assign sub_907_2_n_20 = ~(sub_907_2_n_34 | ~sub_907_2_n_90);
 assign in1_103_9_ = (sub_907_2_n_145 ^ sub_907_2_n_9);
 assign in1_103_17_ = (sub_907_2_n_159 ^ sub_907_2_n_16);
 assign sub_907_2_n_17 = (sub_907_2_n_81 | sub_907_2_n_60);
 assign sub_907_2_n_16 = ~(sub_907_2_n_1 | ~sub_907_2_n_79);
 assign sub_907_2_n_15 = (sub_907_2_n_75 | sub_907_2_n_66);
 assign sub_907_2_n_14 = ~(sub_907_2_n_48 | ~sub_907_2_n_74);
 assign sub_907_2_n_13 = ~(sub_907_2_n_68 | ~sub_907_2_n_69);
 assign sub_907_2_n_12 = ~(sub_907_2_n_61 | ~sub_907_2_n_67);
 assign sub_907_2_n_11 = ~(sub_907_2_n_70 | ~sub_907_2_n_63);
 assign sub_907_2_n_10 = (sub_907_2_n_59 & sub_907_2_n_2);
 assign sub_907_2_n_9 = ~(sub_907_2_n_0 | ~sub_907_2_n_58);
 assign sub_907_2_n_8 = ~(sub_907_2_n_45 | ~sub_907_2_n_55);
 assign sub_907_2_n_7 = ~(sub_907_2_n_66 | ~sub_907_2_n_47);
 assign sub_907_2_n_6 = ~(sub_907_2_n_44 | ~sub_907_2_n_46);
 assign sub_907_2_n_5 = ~(sub_907_2_n_41 | ~sub_907_2_n_42);
 assign sub_907_2_n_4 = ~(sub_907_2_n_50 | ~sub_907_2_n_40);
 assign sub_907_2_n_3 = ~(in1_101_15_ | ~n_1549);
 assign sub_907_2_n_2 = ~(n_1569 & ~in1_101_4_);
 assign sub_907_2_n_1 = ~(in1_101_16_ | ~n_1562);
 assign sub_907_2_n_0 = ~(in1_101_8_ | ~n_1589);
 assign sub_928_2_n_171 = ~(sub_928_2_n_53 & (sub_928_2_n_170 | sub_928_2_n_0));
 assign sub_928_2_n_170 = ~(sub_928_2_n_114 | (sub_928_2_n_164 & sub_928_2_n_100));
 assign sub_928_2_n_169 = ~(sub_928_2_n_52 & ~(sub_928_2_n_164 & sub_928_2_n_82));
 assign sub_928_2_n_168 = ~(sub_928_2_n_64 & (sub_928_2_n_163 | sub_928_2_n_78));
 assign sub_928_2_n_167 = ~(sub_928_2_n_85 & (sub_928_2_n_161 | sub_928_2_n_71));
 assign in1_106_14_ = (sub_928_2_n_161 ^ sub_928_2_n_16);
 assign in1_106_24_ = (sub_928_2_n_157 ^ in1_104_23_);
 assign sub_928_2_n_164 = ~(sub_928_2_n_131 & (sub_928_2_n_42 | sub_928_2_n_120));
 assign sub_928_2_n_163 = ~(sub_928_2_n_113 | ~(sub_928_2_n_42 | sub_928_2_n_96));
 assign sub_928_2_n_162 = ~(sub_928_2_n_51 & (sub_928_2_n_42 | sub_928_2_n_55));
 assign sub_928_2_n_161 = ~(sub_928_2_n_115 | (sub_928_2_n_154 & sub_928_2_n_102));
 assign sub_928_2_n_160 = ~(sub_928_2_n_81 & ~(sub_928_2_n_154 & sub_928_2_n_76));
 assign sub_928_2_n_159 = ~(sub_928_2_n_77 & (sub_928_2_n_40 | sub_928_2_n_56));
 assign in1_106_16_ = ~(sub_928_2_n_42 ^ sub_928_2_n_6);
 assign sub_928_2_n_157 = ~(sub_928_2_n_143 | sub_928_2_n_155);
 assign in1_106_7_ = (sub_928_2_n_152 ^ sub_928_2_n_92);
 assign sub_928_2_n_155 = ~(sub_928_2_n_151 | sub_928_2_n_125);
 assign sub_928_2_n_154 = ~(sub_928_2_n_134 & (sub_928_2_n_149 | sub_928_2_n_29));
 assign sub_928_2_n_153 = ~(sub_928_2_n_57 & (sub_928_2_n_149 | sub_928_2_n_80));
 assign sub_928_2_n_152 = ~(sub_928_2_n_79 & (sub_928_2_n_147 | sub_928_2_n_83));
 assign sub_928_2_n_151 = ~(sub_928_2_n_150 & sub_928_2_n_127);
 assign sub_928_2_n_149 = ~sub_928_2_n_150;
 assign sub_928_2_n_150 = ~(sub_928_2_n_148 & sub_928_2_n_133);
 assign sub_928_2_n_148 = ~(sub_928_2_n_144 & sub_928_2_n_107);
 assign sub_928_2_n_147 = ~(sub_928_2_n_144 | sub_928_2_n_116);
 assign sub_928_2_n_146 = ~(sub_928_2_n_75 | (sub_928_2_n_138 & sub_928_2_n_61));
 assign in1_106_3_ = (sub_928_2_n_141 ^ sub_928_2_n_93);
 assign sub_928_2_n_144 = ~(sub_928_2_n_139 | sub_928_2_n_99);
 assign sub_928_2_n_143 = ~(sub_928_2_n_142 & sub_928_2_n_135);
 assign sub_928_2_n_142 = ~(sub_928_2_n_136 & ~sub_928_2_n_125);
 assign sub_928_2_n_141 = ~(sub_928_2_n_50 & (sub_928_2_n_129 | sub_928_2_n_59));
 assign in1_106_2_ = ~(sub_928_2_n_129 ^ sub_928_2_n_5);
 assign sub_928_2_n_138 = ~sub_928_2_n_139;
 assign sub_928_2_n_139 = ~(sub_928_2_n_137 | sub_928_2_n_110);
 assign sub_928_2_n_137 = ~(sub_928_2_n_129 | sub_928_2_n_12);
 assign sub_928_2_n_136 = ~(sub_928_2_n_132 & (sub_928_2_n_134 | sub_928_2_n_122));
 assign sub_928_2_n_135 = ~(sub_928_2_n_41 | sub_928_2_n_130);
 assign sub_928_2_n_134 = ~(sub_928_2_n_126 | sub_928_2_n_111);
 assign sub_928_2_n_133 = ~(sub_928_2_n_118 | (sub_928_2_n_116 & sub_928_2_n_107));
 assign sub_928_2_n_132 = ~(sub_928_2_n_119 | (sub_928_2_n_115 & sub_928_2_n_105));
 assign sub_928_2_n_131 = ~(sub_928_2_n_117 | (sub_928_2_n_113 & sub_928_2_n_103));
 assign sub_928_2_n_130 = ~(sub_928_2_n_109 & ~(sub_928_2_n_114 & sub_928_2_n_104));
 assign sub_928_2_n_129 = ~(sub_928_2_n_124 | sub_928_2_n_48);
 assign in1_106_1_ = ~(in1_104_0_ ^ (n_1586 ^ sub_928_2_n_49));
 assign sub_928_2_n_127 = ~(sub_928_2_n_29 | sub_928_2_n_122);
 assign sub_928_2_n_126 = ~(sub_928_2_n_112 | sub_928_2_n_11);
 assign sub_928_2_n_125 = ~(sub_928_2_n_121 & ~sub_928_2_n_120);
 assign sub_928_2_n_124 = ~(sub_928_2_n_123 | ~(in1_104_0_ | sub_928_2_n_47));
 assign sub_928_2_n_123 = ~sub_928_2_n_49;
 assign sub_928_2_n_119 = ~(sub_928_2_n_67 & (sub_928_2_n_85 | sub_928_2_n_60));
 assign sub_928_2_n_118 = ~(sub_928_2_n_68 & (sub_928_2_n_79 | sub_928_2_n_70));
 assign sub_928_2_n_117 = ~(sub_928_2_n_90 & (sub_928_2_n_64 | sub_928_2_n_58));
 assign sub_928_2_n_122 = ~(sub_928_2_n_102 & sub_928_2_n_105);
 assign sub_928_2_n_121 = (sub_928_2_n_100 & sub_928_2_n_104);
 assign sub_928_2_n_120 = ~(sub_928_2_n_95 & sub_928_2_n_103);
 assign sub_928_2_n_111 = ~(sub_928_2_n_89 & (sub_928_2_n_77 | sub_928_2_n_1));
 assign sub_928_2_n_110 = ~(sub_928_2_n_91 & (sub_928_2_n_50 | sub_928_2_n_63));
 assign sub_928_2_n_109 = ~(sub_928_2_n_66 | ~(sub_928_2_n_53 | sub_928_2_n_84));
 assign sub_928_2_n_116 = ~(sub_928_2_n_65 & (sub_928_2_n_74 | sub_928_2_n_62));
 assign sub_928_2_n_115 = ~(sub_928_2_n_88 & (sub_928_2_n_81 | sub_928_2_n_54));
 assign sub_928_2_n_114 = ~(sub_928_2_n_69 & (sub_928_2_n_52 | sub_928_2_n_72));
 assign sub_928_2_n_113 = ~(sub_928_2_n_86 & (sub_928_2_n_51 | sub_928_2_n_73));
 assign sub_928_2_n_112 = ~(sub_928_2_n_87 | ~(sub_928_2_n_57 | sub_928_2_n_4));
 assign sub_928_2_n_99 = ~(sub_928_2_n_61 & ~sub_928_2_n_62);
 assign sub_928_2_n_108 = ~(sub_928_2_n_66 | sub_928_2_n_84);
 assign sub_928_2_n_107 = ~(sub_928_2_n_83 | sub_928_2_n_70);
 assign sub_928_2_n_106 = ~(sub_928_2_n_87 | sub_928_2_n_4);
 assign sub_928_2_n_105 = ~(sub_928_2_n_71 | sub_928_2_n_60);
 assign sub_928_2_n_104 = ~(sub_928_2_n_0 | sub_928_2_n_84);
 assign sub_928_2_n_103 = ~(sub_928_2_n_78 | sub_928_2_n_58);
 assign sub_928_2_n_102 = ~(sub_928_2_n_3 | sub_928_2_n_54);
 assign sub_928_2_n_101 = ~(sub_928_2_n_58 | ~sub_928_2_n_90);
 assign sub_928_2_n_100 = ~(sub_928_2_n_2 | sub_928_2_n_72);
 assign sub_928_2_n_96 = ~sub_928_2_n_95;
 assign in1_106_0_ = ~(sub_928_2_n_49 & ~(sub_928_2_n_46 & n_1537));
 assign sub_928_2_n_98 = ~(sub_928_2_n_80 | sub_928_2_n_4);
 assign sub_928_2_n_93 = ~(sub_928_2_n_63 | ~sub_928_2_n_91);
 assign sub_928_2_n_97 = ~(sub_928_2_n_60 | ~sub_928_2_n_67);
 assign sub_928_2_n_92 = ~(sub_928_2_n_70 | ~sub_928_2_n_68);
 assign sub_928_2_n_95 = ~(sub_928_2_n_55 | sub_928_2_n_73);
 assign sub_928_2_n_82 = ~sub_928_2_n_2;
 assign sub_928_2_n_76 = ~sub_928_2_n_3;
 assign sub_928_2_n_75 = ~sub_928_2_n_74;
 assign sub_928_2_n_91 = ~(in1_104_2_ & ~n_1579);
 assign sub_928_2_n_90 = ~(in1_104_18_ & ~n_1558);
 assign sub_928_2_n_89 = ~(in1_104_10_ & ~n_1555);
 assign sub_928_2_n_88 = ~(in1_104_12_ & ~n_1581);
 assign sub_928_2_n_87 = ~(n_1589 | ~in1_104_8_);
 assign sub_928_2_n_86 = ~(in1_104_16_ & ~n_1562);
 assign sub_928_2_n_85 = ~(in1_104_13_ & ~n_1577);
 assign sub_928_2_n_84 = ~(in1_104_22_ | sub_928_2_n_45);
 assign sub_928_2_n_83 = ~(in1_104_5_ | ~n_1567);
 assign sub_928_2_n_81 = ~(in1_104_11_ & ~n_1595);
 assign sub_928_2_n_80 = ~(in1_104_7_ | ~n_1479);
 assign sub_928_2_n_79 = ~(in1_104_5_ & ~n_1567);
 assign sub_928_2_n_78 = ~(in1_104_17_ | ~n_1472);
 assign sub_928_2_n_77 = ~(in1_104_9_ & ~n_1551);
 assign sub_928_2_n_74 = ~(in1_104_3_ & ~n_1535);
 assign sub_928_2_n_73 = ~(in1_104_16_ | ~n_1562);
 assign sub_928_2_n_72 = ~(in1_104_20_ | ~n_1593);
 assign sub_928_2_n_71 = ~(in1_104_13_ | ~n_1577);
 assign sub_928_2_n_70 = ~(in1_104_6_ | ~n_1527);
 assign sub_928_2_n_69 = ~(in1_104_20_ & ~n_1593);
 assign sub_928_2_n_48 = ~(n_1586 | ~in1_104_0_);
 assign sub_928_2_n_68 = ~(in1_104_6_ & ~n_1527);
 assign sub_928_2_n_67 = ~(in1_104_14_ & ~n_1495);
 assign sub_928_2_n_66 = (sub_928_2_n_45 & in1_104_22_);
 assign sub_928_2_n_65 = ~(in1_104_4_ & ~n_1569);
 assign sub_928_2_n_64 = ~(in1_104_17_ & ~n_1472);
 assign sub_928_2_n_63 = ~(in1_104_2_ | ~n_1579);
 assign sub_928_2_n_62 = ~(in1_104_4_ | ~n_1569);
 assign sub_928_2_n_61 = ~(n_1535 & ~in1_104_3_);
 assign sub_928_2_n_60 = ~(in1_104_14_ | ~n_1495);
 assign sub_928_2_n_59 = ~(in1_104_1_ | ~n_1477);
 assign sub_928_2_n_58 = ~(in1_104_18_ | ~n_1558);
 assign sub_928_2_n_57 = ~(in1_104_7_ & ~n_1479);
 assign sub_928_2_n_56 = ~(in1_104_9_ | ~n_1551);
 assign sub_928_2_n_55 = ~(in1_104_15_ | ~n_1549);
 assign sub_928_2_n_54 = ~(in1_104_12_ | ~n_1581);
 assign sub_928_2_n_53 = ~(in1_104_21_ & ~n_1591);
 assign sub_928_2_n_52 = ~(in1_104_19_ & ~n_1565);
 assign sub_928_2_n_51 = ~(in1_104_15_ & ~n_1549);
 assign sub_928_2_n_50 = ~(in1_104_1_ & ~n_1477);
 assign sub_928_2_n_49 = ~(n_1543 & ~n_1537);
 assign sub_928_2_n_47 = ~n_1586;
 assign sub_928_2_n_46 = ~n_1543;
 assign sub_928_2_n_45 = ~n_1403;
 assign in1_106_18_ = ~(sub_928_2_n_163 ^ sub_928_2_n_13);
 assign in1_106_10_ = ~(sub_928_2_n_40 ^ sub_928_2_n_17);
 assign sub_928_2_n_42 = ~(sub_928_2_n_136 | ~sub_928_2_n_151);
 assign sub_928_2_n_41 = ~(sub_928_2_n_131 | ~sub_928_2_n_121);
 assign sub_928_2_n_40 = ~(sub_928_2_n_28 | ~sub_928_2_n_112);
 assign in1_106_8_ = (sub_928_2_n_150 ^ sub_928_2_n_9);
 assign in1_106_23_ = (sub_928_2_n_171 ^ sub_928_2_n_108);
 assign in1_106_9_ = (sub_928_2_n_153 ^ sub_928_2_n_106);
 assign in1_106_6_ = ~(sub_928_2_n_147 ^ sub_928_2_n_18);
 assign in1_106_22_ = ~(sub_928_2_n_170 ^ sub_928_2_n_8);
 assign in1_106_21_ = (sub_928_2_n_169 ^ sub_928_2_n_15);
 assign in1_106_20_ = (sub_928_2_n_164 ^ sub_928_2_n_7);
 assign in1_106_19_ = (sub_928_2_n_168 ^ sub_928_2_n_101);
 assign in1_106_17_ = (sub_928_2_n_162 ^ sub_928_2_n_20);
 assign in1_106_11_ = (sub_928_2_n_159 ^ sub_928_2_n_22);
 assign sub_928_2_n_29 = ~(sub_928_2_n_98 & ~sub_928_2_n_11);
 assign sub_928_2_n_28 = ~(sub_928_2_n_149 | ~sub_928_2_n_98);
 assign in1_106_15_ = (sub_928_2_n_167 ^ sub_928_2_n_97);
 assign in1_106_13_ = (sub_928_2_n_160 ^ sub_928_2_n_21);
 assign in1_106_5_ = ~(sub_928_2_n_146 ^ sub_928_2_n_14);
 assign in1_106_12_ = (sub_928_2_n_154 ^ sub_928_2_n_19);
 assign in1_106_4_ = ~(sub_928_2_n_139 ^ sub_928_2_n_10);
 assign sub_928_2_n_22 = ~(sub_928_2_n_1 | ~sub_928_2_n_89);
 assign sub_928_2_n_21 = ~(sub_928_2_n_54 | ~sub_928_2_n_88);
 assign sub_928_2_n_20 = ~(sub_928_2_n_73 | ~sub_928_2_n_86);
 assign sub_928_2_n_19 = ~(sub_928_2_n_3 | ~sub_928_2_n_81);
 assign sub_928_2_n_18 = ~(sub_928_2_n_83 | ~sub_928_2_n_79);
 assign sub_928_2_n_17 = ~(sub_928_2_n_56 | ~sub_928_2_n_77);
 assign sub_928_2_n_16 = ~(sub_928_2_n_85 & ~sub_928_2_n_71);
 assign sub_928_2_n_15 = ~(sub_928_2_n_72 | ~sub_928_2_n_69);
 assign sub_928_2_n_14 = ~(sub_928_2_n_62 | ~sub_928_2_n_65);
 assign sub_928_2_n_13 = ~(sub_928_2_n_78 | ~sub_928_2_n_64);
 assign sub_928_2_n_12 = (sub_928_2_n_63 | sub_928_2_n_59);
 assign sub_928_2_n_11 = (sub_928_2_n_1 | sub_928_2_n_56);
 assign sub_928_2_n_10 = ~(sub_928_2_n_75 | ~sub_928_2_n_61);
 assign sub_928_2_n_9 = ~(sub_928_2_n_80 | ~sub_928_2_n_57);
 assign sub_928_2_n_8 = ~(sub_928_2_n_0 | ~sub_928_2_n_53);
 assign sub_928_2_n_7 = ~(sub_928_2_n_2 | ~sub_928_2_n_52);
 assign sub_928_2_n_6 = ~(sub_928_2_n_55 | ~sub_928_2_n_51);
 assign sub_928_2_n_5 = ~(sub_928_2_n_59 | ~sub_928_2_n_50);
 assign sub_928_2_n_4 = ~(in1_104_8_ | ~n_1589);
 assign sub_928_2_n_3 = ~(in1_104_11_ | ~n_1595);
 assign sub_928_2_n_2 = ~(in1_104_19_ | ~n_1565);
 assign sub_928_2_n_1 = ~(in1_104_10_ | ~n_1555);
 assign sub_928_2_n_0 = ~(in1_104_21_ | ~n_1591);
 assign sub_949_2_n_170 = ~(sub_949_2_n_62 | (sub_949_2_n_168 & sub_949_2_n_0));
 assign in1_109_21_ = ~(sub_949_2_n_166 ^ sub_949_2_n_19);
 assign in1_109_24_ = ~(sub_949_2_n_160 ^ n_1459);
 assign sub_949_2_n_166 = ~(sub_949_2_n_81 & (sub_949_2_n_161 | sub_949_2_n_77));
 assign sub_949_2_n_165 = ~(n_1447 & (sub_949_2_n_163 | n_1446));
 assign sub_949_2_n_164 = ~(sub_949_2_n_54 & (sub_949_2_n_162 | sub_949_2_n_58));
 assign sub_949_2_n_168 = ~(sub_949_2_n_111 & (sub_949_2_n_161 | sub_949_2_n_91));
 assign sub_949_2_n_160 = ~(sub_949_2_n_152 & sub_949_2_n_140);
 assign sub_949_2_n_159 = ~(n_1453 & (sub_949_2_n_151 | sub_949_2_n_79));
 assign sub_949_2_n_163 = ~(sub_949_2_n_35 | sub_949_2_n_112);
 assign sub_949_2_n_162 = ~(sub_949_2_n_154 | sub_949_2_n_113);
 assign sub_949_2_n_161 = ~(sub_949_2_n_155 | sub_949_2_n_128);
 assign in1_109_16_ = ~(sub_949_2_n_151 ^ sub_949_2_n_5);
 assign sub_949_2_n_157 = ~(sub_949_2_n_57 & (sub_949_2_n_150 | sub_949_2_n_70));
 assign sub_949_2_n_156 = ~(sub_949_2_n_72 & (sub_949_2_n_149 | sub_949_2_n_75));
 assign sub_949_2_n_155 = ~(sub_949_2_n_151 | sub_949_2_n_117);
 assign sub_949_2_n_154 = ~(sub_949_2_n_150 | sub_949_2_n_15);
 assign in1_109_7_ = (sub_949_2_n_146 ^ sub_949_2_n_96);
 assign sub_949_2_n_152 = ~(sub_949_2_n_134 | (n_1424 & sub_949_2_n_37));
 assign sub_949_2_n_151 = ~(n_1424 | n_1417);
 assign sub_949_2_n_150 = ~(sub_949_2_n_36 | sub_949_2_n_127);
 assign sub_949_2_n_149 = ~(sub_949_2_n_22 | sub_949_2_n_119);
 assign sub_949_2_n_148 = ~(sub_949_2_n_83 & (sub_949_2_n_144 | sub_949_2_n_56));
 assign sub_949_2_n_147 = ~(sub_949_2_n_144 | sub_949_2_n_123);
 assign sub_949_2_n_146 = ~(sub_949_2_n_71 & (sub_949_2_n_38 | sub_949_2_n_52));
 assign in1_109_5_ = ~(sub_949_2_n_142 ^ sub_949_2_n_97);
 assign sub_949_2_n_144 = ~(sub_949_2_n_143 | sub_949_2_n_126);
 assign sub_949_2_n_143 = ~(sub_949_2_n_141 | sub_949_2_n_4);
 assign sub_949_2_n_142 = ~(sub_949_2_n_45 & (sub_949_2_n_138 | sub_949_2_n_47));
 assign sub_949_2_n_141 = ~(sub_949_2_n_137 & sub_949_2_n_98);
 assign sub_949_2_n_140 = ~(n_1417 & sub_949_2_n_37);
 assign sub_949_2_n_139 = ~(sub_949_2_n_60 | (sub_949_2_n_133 & sub_949_2_n_74));
 assign sub_949_2_n_138 = ~sub_949_2_n_137;
 assign sub_949_2_n_137 = ~(sub_949_2_n_135 & sub_949_2_n_116);
 assign sub_949_2_n_136 = ~(sub_949_2_n_130 & ~(sub_949_2_n_127 & sub_949_2_n_121));
 assign sub_949_2_n_135 = ~(sub_949_2_n_133 & sub_949_2_n_99);
 assign sub_949_2_n_134 = ~(sub_949_2_n_129 & ~(sub_949_2_n_128 & sub_949_2_n_120));
 assign sub_949_2_n_133 = ~(sub_949_2_n_132 & sub_949_2_n_44);
 assign sub_949_2_n_132 = ~(sub_949_2_n_125 | (sub_949_2_n_68 & in1_107_0_));
 assign in1_109_1_ = ~(n_1467 ^ (n_1587 ^ n_1540));
 assign sub_949_2_n_130 = ~(sub_949_2_n_107 | (sub_949_2_n_113 & sub_949_2_n_95));
 assign sub_949_2_n_129 = ~(sub_949_2_n_124 | sub_949_2_n_109);
 assign sub_949_2_n_128 = ~(sub_949_2_n_110 & ~(sub_949_2_n_112 & sub_949_2_n_101));
 assign sub_949_2_n_127 = ~(sub_949_2_n_115 & ~(sub_949_2_n_119 & sub_949_2_n_103));
 assign sub_949_2_n_126 = ~(sub_949_2_n_122 & sub_949_2_n_108);
 assign sub_949_2_n_125 = ~(n_1586 | ~sub_949_2_n_68);
 assign sub_949_2_n_124 = ~(sub_949_2_n_111 | sub_949_2_n_102);
 assign sub_949_2_n_123 = ~(sub_949_2_n_118 & sub_949_2_n_121);
 assign sub_949_2_n_122 = ~(sub_949_2_n_114 & ~sub_949_2_n_4);
 assign sub_949_2_n_116 = ~(sub_949_2_n_85 | ~(sub_949_2_n_59 | sub_949_2_n_1));
 assign sub_949_2_n_115 = ~(sub_949_2_n_88 | ~(sub_949_2_n_72 | sub_949_2_n_46));
 assign sub_949_2_n_121 = ~(sub_949_2_n_15 | ~sub_949_2_n_95);
 assign sub_949_2_n_120 = ~(sub_949_2_n_91 | sub_949_2_n_102);
 assign sub_949_2_n_119 = ~(sub_949_2_n_84 & (sub_949_2_n_83 | sub_949_2_n_69));
 assign sub_949_2_n_118 = (sub_949_2_n_93 & sub_949_2_n_103);
 assign sub_949_2_n_117 = ~(sub_949_2_n_106 & sub_949_2_n_101);
 assign sub_949_2_n_110 = ~(sub_949_2_n_67 | ~(n_1447 | n_1466));
 assign sub_949_2_n_109 = ~(sub_949_2_n_64 & (sub_949_2_n_61 | n_1405));
 assign sub_949_2_n_108 = ~(sub_949_2_n_86 | ~(sub_949_2_n_71 | sub_949_2_n_48));
 assign sub_949_2_n_107 = ~(sub_949_2_n_65 & (sub_949_2_n_54 | sub_949_2_n_78));
 assign sub_949_2_n_114 = ~(sub_949_2_n_66 & (sub_949_2_n_45 | sub_949_2_n_2));
 assign sub_949_2_n_113 = ~(sub_949_2_n_89 & (sub_949_2_n_57 | sub_949_2_n_80));
 assign sub_949_2_n_112 = ~(n_1457 & (n_1453 | n_1458));
 assign sub_949_2_n_111 = ~(sub_949_2_n_87 | ~(sub_949_2_n_81 | sub_949_2_n_53));
 assign sub_949_2_n_99 = ~(sub_949_2_n_73 | sub_949_2_n_1);
 assign sub_949_2_n_98 = ~(sub_949_2_n_47 | sub_949_2_n_2);
 assign sub_949_2_n_106 = ~(sub_949_2_n_79 | n_1458);
 assign sub_949_2_n_105 = ~(sub_949_2_n_85 | sub_949_2_n_1);
 assign sub_949_2_n_97 = ~(sub_949_2_n_66 & ~sub_949_2_n_2);
 assign sub_949_2_n_104 = ~(sub_949_2_n_60 | sub_949_2_n_73);
 assign sub_949_2_n_103 = ~(sub_949_2_n_75 | sub_949_2_n_46);
 assign sub_949_2_n_102 = ~(sub_949_2_n_0 & ~n_1405);
 assign sub_949_2_n_96 = ~(sub_949_2_n_86 | sub_949_2_n_48);
 assign sub_949_2_n_101 = ~(n_1446 | n_1466);
 assign sub_949_2_n_100 = ~(sub_949_2_n_67 | n_1466);
 assign in1_109_0_ = ~(n_1540 & ~(sub_949_2_n_43 & n_1539));
 assign sub_949_2_n_95 = ~(sub_949_2_n_58 | sub_949_2_n_78);
 assign sub_949_2_n_94 = ~(sub_949_2_n_88 | sub_949_2_n_46);
 assign sub_949_2_n_93 = ~(sub_949_2_n_56 | sub_949_2_n_69);
 assign sub_949_2_n_92 = ~(sub_949_2_n_80 | ~sub_949_2_n_89);
 assign sub_949_2_n_91 = (sub_949_2_n_77 | sub_949_2_n_53);
 assign sub_949_2_n_74 = ~sub_949_2_n_73;
 assign sub_949_2_n_89 = ~(in1_107_12_ & ~n_1581);
 assign sub_949_2_n_88 = ~(n_1555 | ~in1_107_10_);
 assign sub_949_2_n_87 = ~(n_1594 | ~n_1444);
 assign sub_949_2_n_86 = ~(n_1527 | ~in1_107_6_);
 assign sub_949_2_n_85 = ~(n_1579 | ~in1_107_2_);
 assign sub_949_2_n_84 = ~(in1_107_8_ & ~n_1589);
 assign sub_949_2_n_83 = ~(in1_107_7_ & ~n_1479);
 assign sub_949_2_n_82 = ~(in1_107_18_ | ~n_1558);
 assign sub_949_2_n_81 = ~(n_1450 & ~n_1566);
 assign sub_949_2_n_80 = ~(in1_107_12_ | ~n_1581);
 assign sub_949_2_n_79 = ~(n_1421 | ~n_1550);
 assign sub_949_2_n_78 = ~(in1_107_14_ | ~n_1495);
 assign sub_949_2_n_77 = ~(n_1450 | ~n_1566);
 assign sub_949_2_n_76 = ~(in1_107_22_ | ~n_1403);
 assign sub_949_2_n_75 = ~(in1_107_9_ | ~n_1551);
 assign sub_949_2_n_73 = ~(in1_107_1_ | ~n_1477);
 assign sub_949_2_n_72 = ~(in1_107_9_ & ~n_1551);
 assign sub_949_2_n_71 = ~(in1_107_5_ & ~n_1567);
 assign sub_949_2_n_70 = ~(in1_107_11_ | ~n_1595);
 assign sub_949_2_n_69 = ~(in1_107_8_ | ~n_1589);
 assign sub_949_2_n_68 = ~(n_1543 & ~n_1538);
 assign sub_949_2_n_62 = ~sub_949_2_n_61;
 assign sub_949_2_n_60 = ~sub_949_2_n_59;
 assign sub_949_2_n_44 = ~(in1_107_0_ & ~n_1586);
 assign sub_949_2_n_67 = ~(n_1559 | ~n_1441);
 assign sub_949_2_n_66 = ~(in1_107_4_ & ~n_1569);
 assign sub_949_2_n_65 = ~(in1_107_14_ & ~n_1495);
 assign sub_949_2_n_64 = ~(n_1439 & ~n_1404);
 assign sub_949_2_n_63 = ~(in1_107_16_ & ~n_1562);
 assign sub_949_2_n_61 = ~(n_1442 & ~n_1592);
 assign sub_949_2_n_59 = ~(in1_107_1_ & ~n_1477);
 assign sub_949_2_n_58 = ~(in1_107_13_ | ~n_1577);
 assign sub_949_2_n_57 = ~(in1_107_11_ & ~n_1595);
 assign sub_949_2_n_56 = ~(in1_107_7_ | ~n_1479);
 assign sub_949_2_n_55 = ~(in1_107_16_ | ~n_1562);
 assign sub_949_2_n_54 = ~(in1_107_13_ & ~n_1577);
 assign sub_949_2_n_53 = ~(n_1444 | ~n_1594);
 assign sub_949_2_n_52 = ~(in1_107_5_ | ~n_1567);
 assign sub_949_2_n_51 = ~(in1_107_17_ & ~n_1472);
 assign sub_949_2_n_50 = ~(in1_107_17_ | ~n_1472);
 assign sub_949_2_n_49 = ~(in1_107_15_ & ~n_1549);
 assign sub_949_2_n_48 = ~(in1_107_6_ | ~n_1527);
 assign sub_949_2_n_47 = ~(in1_107_3_ | ~n_1535);
 assign sub_949_2_n_46 = ~(in1_107_10_ | ~n_1555);
 assign sub_949_2_n_45 = ~(in1_107_3_ & ~n_1535);
 assign sub_949_2_n_43 = ~n_1544;
 assign in1_109_18_ = ~(sub_949_2_n_163 ^ sub_949_2_n_6);
 assign in1_109_12_ = ~(sub_949_2_n_150 ^ sub_949_2_n_8);
 assign in1_109_10_ = ~(sub_949_2_n_149 ^ sub_949_2_n_14);
 assign in1_109_8_ = ~(sub_949_2_n_144 ^ sub_949_2_n_17);
 assign sub_949_2_n_38 = ~(sub_949_2_n_114 | ~sub_949_2_n_141);
 assign sub_949_2_n_37 = ~(sub_949_2_n_117 | ~sub_949_2_n_120);
 assign sub_949_2_n_36 = ~(sub_949_2_n_144 | ~sub_949_2_n_118);
 assign sub_949_2_n_35 = ~(sub_949_2_n_151 | ~sub_949_2_n_106);
 assign in1_109_6_ = ~(sub_949_2_n_38 ^ sub_949_2_n_13);
 assign in1_109_3_ = ~(sub_949_2_n_139 ^ sub_949_2_n_105);
 assign in1_109_2_ = (sub_949_2_n_133 ^ sub_949_2_n_104);
 assign in1_109_23_ = ~(sub_949_2_n_170 ^ sub_949_2_n_11);
 assign in1_109_9_ = (sub_949_2_n_148 ^ sub_949_2_n_18);
 assign in1_109_22_ = (sub_949_2_n_168 ^ sub_949_2_n_9);
 assign in1_109_20_ = ~(sub_949_2_n_161 ^ sub_949_2_n_16);
 assign in1_109_19_ = (sub_949_2_n_165 ^ sub_949_2_n_100);
 assign in1_109_4_ = ~(sub_949_2_n_138 ^ sub_949_2_n_3);
 assign in1_109_17_ = (sub_949_2_n_159 ^ sub_949_2_n_10);
 assign in1_109_11_ = (sub_949_2_n_156 ^ sub_949_2_n_94);
 assign in1_109_14_ = ~(n_1418 ^ n_1437);
 assign sub_949_2_n_22 = ~(sub_949_2_n_144 | ~sub_949_2_n_93);
 assign in1_109_13_ = (sub_949_2_n_157 ^ sub_949_2_n_92);
 assign in1_109_15_ = (n_1419 ^ n_1423);
 assign sub_949_2_n_19 = (sub_949_2_n_87 | sub_949_2_n_53);
 assign sub_949_2_n_18 = ~(sub_949_2_n_69 | ~sub_949_2_n_84);
 assign sub_949_2_n_17 = ~(sub_949_2_n_56 | ~sub_949_2_n_83);
 assign sub_949_2_n_16 = ~(sub_949_2_n_77 | ~sub_949_2_n_81);
 assign sub_949_2_n_15 = (sub_949_2_n_80 | sub_949_2_n_70);
 assign sub_949_2_n_14 = ~(sub_949_2_n_75 | ~sub_949_2_n_72);
 assign sub_949_2_n_13 = ~(sub_949_2_n_52 | ~sub_949_2_n_71);
 assign sub_949_2_n_12 = ~(sub_949_2_n_78 | ~sub_949_2_n_65);
 assign sub_949_2_n_11 = ~(n_1405 | ~sub_949_2_n_64);
 assign sub_949_2_n_10 = ~(n_1458 | ~n_1457);
 assign sub_949_2_n_9 = ~(sub_949_2_n_62 | ~sub_949_2_n_0);
 assign sub_949_2_n_8 = ~(sub_949_2_n_70 | ~sub_949_2_n_57);
 assign sub_949_2_n_7 = ~(sub_949_2_n_58 | ~sub_949_2_n_54);
 assign sub_949_2_n_6 = ~(n_1446 | ~n_1447);
 assign sub_949_2_n_5 = ~(sub_949_2_n_79 | ~n_1453);
 assign sub_949_2_n_4 = (sub_949_2_n_48 | sub_949_2_n_52);
 assign sub_949_2_n_3 = ~(sub_949_2_n_47 | ~sub_949_2_n_45);
 assign sub_949_2_n_2 = ~(in1_107_4_ | ~n_1569);
 assign sub_949_2_n_1 = ~(in1_107_2_ | ~n_1579);
 assign sub_949_2_n_0 = ~(n_1592 & ~n_1442);
 assign sub_970_2_n_183 = ~(sub_970_2_n_34 | (sub_970_2_n_180 & sub_970_2_n_61));
 assign in1_112_19_ = ~(sub_970_2_n_178 ^ sub_970_2_n_100);
 assign in1_112_15_ = ~(sub_970_2_n_177 ^ sub_970_2_n_86);
 assign sub_970_2_n_180 = ~(sub_970_2_n_120 & (sub_970_2_n_171 | sub_970_2_n_94));
 assign sub_970_2_n_179 = ~(sub_970_2_n_173 | sub_970_2_n_33);
 assign sub_970_2_n_178 = ~(sub_970_2_n_47 | ~(sub_970_2_n_170 | sub_970_2_n_66));
 assign sub_970_2_n_177 = ~(sub_970_2_n_75 & (sub_970_2_n_21 | sub_970_2_n_56));
 assign in1_112_14_ = ~(sub_970_2_n_21 ^ sub_970_2_n_4);
 assign in1_112_13_ = ~(sub_970_2_n_168 ^ sub_970_2_n_85);
 assign in1_112_11_ = ~(sub_970_2_n_167 ^ sub_970_2_n_6);
 assign sub_970_2_n_173 = ~(sub_970_2_n_171 | sub_970_2_n_73);
 assign in1_112_24_ = (sub_970_2_n_161 ^ in1_110_23_);
 assign sub_970_2_n_171 = ~(sub_970_2_n_135 | ~(sub_970_2_n_160 | sub_970_2_n_126));
 assign sub_970_2_n_170 = ~(sub_970_2_n_8 | sub_970_2_n_119);
 assign sub_970_2_n_169 = ~(sub_970_2_n_162 | sub_970_2_n_49);
 assign sub_970_2_n_168 = ~(sub_970_2_n_72 | (sub_970_2_n_159 & sub_970_2_n_63));
 assign sub_970_2_n_167 = ~(sub_970_2_n_65 | (sub_970_2_n_158 & sub_970_2_n_1));
 assign in1_112_16_ = ~(sub_970_2_n_160 ^ sub_970_2_n_99);
 assign in1_112_12_ = ~(sub_970_2_n_159 ^ sub_970_2_n_83);
 assign in1_112_10_ = ~(sub_970_2_n_158 ^ sub_970_2_n_84);
 assign in1_112_9_ = ~(sub_970_2_n_157 ^ sub_970_2_n_101);
 assign sub_970_2_n_162 = ~(sub_970_2_n_160 | sub_970_2_n_37);
 assign sub_970_2_n_161 = ~(sub_970_2_n_146 | (sub_970_2_n_153 & sub_970_2_n_130));
 assign sub_970_2_n_160 = ~(sub_970_2_n_153 | sub_970_2_n_142);
 assign sub_970_2_n_159 = ~sub_970_2_n_22;
 assign sub_970_2_n_158 = ~(sub_970_2_n_118 & (sub_970_2_n_152 | sub_970_2_n_97));
 assign sub_970_2_n_157 = ~(sub_970_2_n_38 & (sub_970_2_n_152 | sub_970_2_n_69));
 assign in1_112_8_ = ~(sub_970_2_n_152 ^ sub_970_2_n_2);
 assign sub_970_2_n_155 = ~(sub_970_2_n_152 | sub_970_2_n_12);
 assign sub_970_2_n_154 = ~(sub_970_2_n_68 | (sub_970_2_n_150 & sub_970_2_n_0));
 assign sub_970_2_n_153 = ~(sub_970_2_n_152 | sub_970_2_n_132);
 assign sub_970_2_n_152 = ~(sub_970_2_n_151 | sub_970_2_n_137);
 assign sub_970_2_n_151 = ~(sub_970_2_n_147 | sub_970_2_n_113);
 assign sub_970_2_n_150 = ~(sub_970_2_n_147 & sub_970_2_n_122);
 assign sub_970_2_n_149 = ~(sub_970_2_n_40 | (sub_970_2_n_144 & sub_970_2_n_44));
 assign in1_112_4_ = ~(sub_970_2_n_144 ^ sub_970_2_n_82);
 assign sub_970_2_n_147 = ~(sub_970_2_n_144 & sub_970_2_n_103);
 assign sub_970_2_n_146 = ~(sub_970_2_n_141 & ~(sub_970_2_n_142 & sub_970_2_n_130));
 assign sub_970_2_n_145 = ~(sub_970_2_n_29 | (sub_970_2_n_140 & sub_970_2_n_36));
 assign sub_970_2_n_144 = ~(sub_970_2_n_143 & sub_970_2_n_116);
 assign sub_970_2_n_143 = ~(sub_970_2_n_140 & sub_970_2_n_89);
 assign sub_970_2_n_142 = ~(sub_970_2_n_136 & (sub_970_2_n_138 | sub_970_2_n_19));
 assign sub_970_2_n_141 = ~(sub_970_2_n_134 | (sub_970_2_n_135 & sub_970_2_n_128));
 assign sub_970_2_n_140 = ((sub_970_2_n_27 & in1_110_0_) | ((in1_110_0_ & sub_970_2_n_26) | (sub_970_2_n_26
    & sub_970_2_n_27)));
 assign in1_112_1_ = (in1_110_0_ ^ (sub_970_2_n_26 ^ sub_970_2_n_27));
 assign sub_970_2_n_138 = ~(sub_970_2_n_131 | sub_970_2_n_117);
 assign sub_970_2_n_137 = ~(sub_970_2_n_124 & (sub_970_2_n_122 | sub_970_2_n_113));
 assign sub_970_2_n_136 = ~(sub_970_2_n_133 | sub_970_2_n_125);
 assign sub_970_2_n_135 = ~(sub_970_2_n_123 & ~(sub_970_2_n_119 & sub_970_2_n_108));
 assign sub_970_2_n_134 = ~(sub_970_2_n_129 & sub_970_2_n_115);
 assign sub_970_2_n_133 = ~(sub_970_2_n_121 | sub_970_2_n_112);
 assign sub_970_2_n_132 = (sub_970_2_n_12 | sub_970_2_n_19);
 assign sub_970_2_n_131 = ~(sub_970_2_n_118 | sub_970_2_n_98);
 assign sub_970_2_n_130 = ~(sub_970_2_n_126 | sub_970_2_n_127);
 assign sub_970_2_n_129 = ~(sub_970_2_n_111 & ~sub_970_2_n_120);
 assign sub_970_2_n_128 = ~sub_970_2_n_127;
 assign sub_970_2_n_125 = ~(sub_970_2_n_53 & (sub_970_2_n_75 | sub_970_2_n_42));
 assign sub_970_2_n_124 = ~(sub_970_2_n_55 | ~(sub_970_2_n_67 | sub_970_2_n_70));
 assign sub_970_2_n_123 = ~(sub_970_2_n_80 | (sub_970_2_n_47 & sub_970_2_n_30));
 assign sub_970_2_n_127 = ~(sub_970_2_n_111 & ~sub_970_2_n_94);
 assign sub_970_2_n_126 = ~(sub_970_2_n_91 & sub_970_2_n_108);
 assign sub_970_2_n_117 = ~(sub_970_2_n_79 & (sub_970_2_n_64 | sub_970_2_n_45));
 assign sub_970_2_n_116 = ~(sub_970_2_n_81 | ~(sub_970_2_n_28 | sub_970_2_n_46));
 assign sub_970_2_n_115 = ~(sub_970_2_n_88 | sub_970_2_n_52);
 assign sub_970_2_n_122 = ~(sub_970_2_n_104 | sub_970_2_n_51);
 assign sub_970_2_n_121 = ~(sub_970_2_n_78 | ~(sub_970_2_n_71 | sub_970_2_n_50));
 assign sub_970_2_n_120 = ~(sub_970_2_n_102 | sub_970_2_n_54);
 assign sub_970_2_n_119 = ~(sub_970_2_n_76 & (sub_970_2_n_48 | sub_970_2_n_58));
 assign sub_970_2_n_118 = ~(sub_970_2_n_77 | ~(sub_970_2_n_38 | sub_970_2_n_59));
 assign sub_970_2_n_104 = ~(sub_970_2_n_39 | sub_970_2_n_41);
 assign sub_970_2_n_103 = ~(sub_970_2_n_43 | sub_970_2_n_41);
 assign sub_970_2_n_102 = ~(sub_970_2_n_32 | sub_970_2_n_57);
 assign sub_970_2_n_114 = ~(sub_970_2_n_34 | sub_970_2_n_60);
 assign sub_970_2_n_113 = ~(sub_970_2_n_0 & ~sub_970_2_n_70);
 assign sub_970_2_n_101 = (sub_970_2_n_77 | sub_970_2_n_59);
 assign sub_970_2_n_112 = (sub_970_2_n_56 | sub_970_2_n_42);
 assign sub_970_2_n_111 = ~(sub_970_2_n_60 | sub_970_2_n_74);
 assign sub_970_2_n_110 = ~(sub_970_2_n_52 | sub_970_2_n_74);
 assign sub_970_2_n_109 = ~(sub_970_2_n_54 | sub_970_2_n_57);
 assign sub_970_2_n_108 = ~(sub_970_2_n_66 | sub_970_2_n_31);
 assign sub_970_2_n_107 = ~(sub_970_2_n_62 | sub_970_2_n_50);
 assign sub_970_2_n_106 = ~(sub_970_2_n_33 | sub_970_2_n_73);
 assign sub_970_2_n_105 = ~(sub_970_2_n_29 | sub_970_2_n_35);
 assign sub_970_2_n_100 = ~(sub_970_2_n_80 | sub_970_2_n_31);
 assign sub_970_2_n_99 = ~(sub_970_2_n_49 | sub_970_2_n_37);
 assign sub_970_2_n_97 = ~sub_970_2_n_96;
 assign sub_970_2_n_89 = ~(sub_970_2_n_35 | sub_970_2_n_46);
 assign sub_970_2_n_88 = ~(sub_970_2_n_74 | ~sub_970_2_n_34);
 assign in1_112_0_ = ~(sub_970_2_n_27 & ~(sub_970_2_n_25 & n_1523));
 assign sub_970_2_n_98 = ~(sub_970_2_n_1 & ~sub_970_2_n_45);
 assign sub_970_2_n_96 = ~(sub_970_2_n_69 | sub_970_2_n_59);
 assign sub_970_2_n_95 = ~(sub_970_2_n_81 | sub_970_2_n_46);
 assign sub_970_2_n_86 = ~(sub_970_2_n_53 & ~sub_970_2_n_42);
 assign sub_970_2_n_94 = (sub_970_2_n_73 | sub_970_2_n_57);
 assign sub_970_2_n_93 = ~(sub_970_2_n_55 | sub_970_2_n_70);
 assign sub_970_2_n_85 = ~(sub_970_2_n_78 | sub_970_2_n_50);
 assign sub_970_2_n_92 = ~(sub_970_2_n_51 | sub_970_2_n_41);
 assign sub_970_2_n_91 = ~(sub_970_2_n_37 | sub_970_2_n_58);
 assign sub_970_2_n_84 = ~(sub_970_2_n_64 & sub_970_2_n_1);
 assign sub_970_2_n_83 = ~(sub_970_2_n_71 & sub_970_2_n_63);
 assign sub_970_2_n_90 = ~(sub_970_2_n_47 | sub_970_2_n_66);
 assign sub_970_2_n_82 = ~(sub_970_2_n_39 & sub_970_2_n_44);
 assign sub_970_2_n_72 = ~sub_970_2_n_71;
 assign sub_970_2_n_68 = ~sub_970_2_n_67;
 assign sub_970_2_n_65 = ~sub_970_2_n_64;
 assign sub_970_2_n_63 = ~sub_970_2_n_62;
 assign sub_970_2_n_61 = ~sub_970_2_n_60;
 assign sub_970_2_n_81 = ~(n_1580 | ~in1_110_2_);
 assign sub_970_2_n_80 = ~(n_1559 | ~in1_110_18_);
 assign sub_970_2_n_79 = ~(in1_110_10_ & ~n_1556);
 assign sub_970_2_n_78 = ~(n_1582 | ~in1_110_12_);
 assign sub_970_2_n_77 = ~(n_1590 | ~in1_110_8_);
 assign sub_970_2_n_76 = ~(in1_110_16_ & ~n_1563);
 assign sub_970_2_n_75 = ~(in1_110_13_ & ~n_1578);
 assign sub_970_2_n_74 = ~(in1_110_22_ | sub_970_2_n_24);
 assign sub_970_2_n_73 = ~(in1_110_19_ | ~n_1566);
 assign sub_970_2_n_71 = ~(in1_110_11_ & ~n_1596);
 assign sub_970_2_n_70 = ~(in1_110_6_ | ~n_1528);
 assign sub_970_2_n_69 = ~(in1_110_7_ | ~n_1480);
 assign sub_970_2_n_67 = ~(in1_110_5_ & ~n_1568);
 assign sub_970_2_n_66 = ~(in1_110_17_ | ~n_1473);
 assign sub_970_2_n_64 = ~(in1_110_9_ & ~n_1552);
 assign sub_970_2_n_62 = ~(in1_110_11_ | ~n_1596);
 assign sub_970_2_n_60 = ~(in1_110_21_ | ~n_1592);
 assign sub_970_2_n_59 = ~(in1_110_8_ | ~n_1590);
 assign sub_970_2_n_58 = ~(in1_110_16_ | ~n_1563);
 assign sub_970_2_n_57 = ~(in1_110_20_ | ~n_1594);
 assign sub_970_2_n_56 = ~(in1_110_13_ | ~n_1578);
 assign sub_970_2_n_49 = ~sub_970_2_n_48;
 assign sub_970_2_n_44 = ~sub_970_2_n_43;
 assign sub_970_2_n_40 = ~sub_970_2_n_39;
 assign sub_970_2_n_36 = ~sub_970_2_n_35;
 assign sub_970_2_n_33 = ~sub_970_2_n_32;
 assign sub_970_2_n_30 = ~sub_970_2_n_31;
 assign sub_970_2_n_29 = ~sub_970_2_n_28;
 assign sub_970_2_n_55 = ~(n_1528 | ~in1_110_6_);
 assign sub_970_2_n_54 = ~(n_1594 | ~in1_110_20_);
 assign sub_970_2_n_53 = ~(in1_110_14_ & ~n_1496);
 assign sub_970_2_n_52 = (sub_970_2_n_24 & in1_110_22_);
 assign sub_970_2_n_51 = ~(n_1570 | ~in1_110_4_);
 assign sub_970_2_n_50 = ~(in1_110_12_ | ~n_1582);
 assign sub_970_2_n_48 = ~(in1_110_15_ & ~n_1550);
 assign sub_970_2_n_47 = ~(n_1473 | ~in1_110_17_);
 assign sub_970_2_n_46 = ~(in1_110_2_ | ~n_1580);
 assign sub_970_2_n_45 = ~(in1_110_10_ | ~n_1556);
 assign sub_970_2_n_43 = ~(in1_110_3_ | ~n_1536);
 assign sub_970_2_n_42 = ~(in1_110_14_ | ~n_1496);
 assign sub_970_2_n_41 = ~(in1_110_4_ | ~n_1570);
 assign sub_970_2_n_39 = ~(in1_110_3_ & ~n_1536);
 assign sub_970_2_n_38 = ~(in1_110_7_ & ~n_1480);
 assign sub_970_2_n_37 = ~(in1_110_15_ | ~n_1550);
 assign sub_970_2_n_35 = ~(in1_110_1_ | ~n_1478);
 assign sub_970_2_n_34 = ~(n_1592 | ~in1_110_21_);
 assign sub_970_2_n_32 = ~(in1_110_19_ & ~n_1566);
 assign sub_970_2_n_31 = ~(in1_110_18_ | ~n_1559);
 assign sub_970_2_n_28 = ~(in1_110_1_ & ~n_1478);
 assign sub_970_2_n_27 = ~(n_1544 & ~n_1523);
 assign sub_970_2_n_26 = ~n_1587;
 assign sub_970_2_n_25 = ~n_1544;
 assign sub_970_2_n_24 = ~n_1404;
 assign in1_112_6_ = (sub_970_2_n_150 ^ sub_970_2_n_3);
 assign sub_970_2_n_22 = ~(sub_970_2_n_155 | ~sub_970_2_n_138);
 assign sub_970_2_n_21 = ~(sub_970_2_n_16 | ~sub_970_2_n_121);
 assign in1_112_22_ = (sub_970_2_n_180 ^ sub_970_2_n_114);
 assign sub_970_2_n_19 = ~(sub_970_2_n_107 & ~sub_970_2_n_112);
 assign in1_112_23_ = ~(sub_970_2_n_183 ^ sub_970_2_n_110);
 assign in1_112_21_ = ~(sub_970_2_n_179 ^ sub_970_2_n_109);
 assign sub_970_2_n_16 = ~(sub_970_2_n_22 | ~sub_970_2_n_107);
 assign in1_112_20_ = ~(sub_970_2_n_171 ^ sub_970_2_n_106);
 assign in1_112_2_ = (sub_970_2_n_140 ^ sub_970_2_n_105);
 assign in1_112_17_ = ~(sub_970_2_n_169 ^ sub_970_2_n_5);
 assign sub_970_2_n_12 = ~(sub_970_2_n_96 & ~sub_970_2_n_98);
 assign in1_112_3_ = ~(sub_970_2_n_145 ^ sub_970_2_n_95);
 assign in1_112_7_ = ~(sub_970_2_n_154 ^ sub_970_2_n_93);
 assign in1_112_5_ = ~(sub_970_2_n_149 ^ sub_970_2_n_92);
 assign sub_970_2_n_8 = ~(sub_970_2_n_160 | ~sub_970_2_n_91);
 assign in1_112_18_ = ~(sub_970_2_n_170 ^ sub_970_2_n_90);
 assign sub_970_2_n_6 = ~(sub_970_2_n_45 | ~sub_970_2_n_79);
 assign sub_970_2_n_5 = ~(sub_970_2_n_58 | ~sub_970_2_n_76);
 assign sub_970_2_n_4 = ~(sub_970_2_n_56 | ~sub_970_2_n_75);
 assign sub_970_2_n_3 = ~(sub_970_2_n_68 | ~sub_970_2_n_0);
 assign sub_970_2_n_2 = ~(sub_970_2_n_69 | ~sub_970_2_n_38);
 assign sub_970_2_n_1 = ~(n_1552 & ~in1_110_9_);
 assign sub_970_2_n_0 = ~(n_1568 & ~in1_110_5_);
 assign sub_991_2_n_172 = ~(sub_991_2_n_56 & (sub_991_2_n_171 | sub_991_2_n_5));
 assign sub_991_2_n_171 = ~(sub_991_2_n_118 | (sub_991_2_n_166 & sub_991_2_n_98));
 assign sub_991_2_n_170 = ~(sub_991_2_n_81 & (sub_991_2_n_165 | sub_991_2_n_3));
 assign sub_991_2_n_169 = ~(sub_991_2_n_75 & (sub_991_2_n_164 | sub_991_2_n_54));
 assign in1_115_24_ = ~(sub_991_2_n_161 ^ in1_113_23_);
 assign sub_991_2_n_167 = ~(sub_991_2_n_57 & (sub_991_2_n_159 | sub_991_2_n_2));
 assign sub_991_2_n_165 = ~sub_991_2_n_166;
 assign sub_991_2_n_166 = ~(sub_991_2_n_130 & (sub_991_2_n_156 | sub_991_2_n_32));
 assign sub_991_2_n_164 = ~sub_991_2_n_163;
 assign sub_991_2_n_163 = ~(sub_991_2_n_115 & (sub_991_2_n_156 | sub_991_2_n_96));
 assign sub_991_2_n_162 = ~(sub_991_2_n_55 & (sub_991_2_n_156 | sub_991_2_n_82));
 assign sub_991_2_n_161 = ~(sub_991_2_n_155 & (sub_991_2_n_138 & sub_991_2_n_144));
 assign in1_115_16_ = ~(sub_991_2_n_156 ^ sub_991_2_n_9);
 assign sub_991_2_n_159 = ~(sub_991_2_n_25 | sub_991_2_n_116);
 assign sub_991_2_n_158 = ~(sub_991_2_n_52 & (sub_991_2_n_44 | sub_991_2_n_50));
 assign sub_991_2_n_157 = ~(sub_991_2_n_86 | (sub_991_2_n_153 & sub_991_2_n_1));
 assign sub_991_2_n_156 = ~(sub_991_2_n_154 | sub_991_2_n_140);
 assign sub_991_2_n_155 = ~(sub_991_2_n_154 & sub_991_2_n_125);
 assign sub_991_2_n_154 = ~(sub_991_2_n_151 | sub_991_2_n_122);
 assign sub_991_2_n_153 = ~(sub_991_2_n_124 & (sub_991_2_n_147 | sub_991_2_n_97));
 assign sub_991_2_n_152 = ~(sub_991_2_n_53 & (sub_991_2_n_147 | sub_991_2_n_70));
 assign sub_991_2_n_151 = ~(sub_991_2_n_148 & sub_991_2_n_120);
 assign sub_991_2_n_150 = ~(sub_991_2_n_60 & (sub_991_2_n_43 | sub_991_2_n_80));
 assign in1_115_5_ = ~(sub_991_2_n_146 ^ sub_991_2_n_91);
 assign sub_991_2_n_147 = ~sub_991_2_n_148;
 assign sub_991_2_n_148 = ~(sub_991_2_n_129 & (sub_991_2_n_145 | sub_991_2_n_10));
 assign sub_991_2_n_146 = ~(sub_991_2_n_71 & (sub_991_2_n_142 | sub_991_2_n_84));
 assign sub_991_2_n_145 = ~(sub_991_2_n_141 & sub_991_2_n_102);
 assign sub_991_2_n_144 = ~(sub_991_2_n_140 & sub_991_2_n_125);
 assign sub_991_2_n_143 = ~(sub_991_2_n_78 | (sub_991_2_n_136 & sub_991_2_n_73));
 assign sub_991_2_n_142 = ~sub_991_2_n_141;
 assign sub_991_2_n_141 = ~(sub_991_2_n_139 & sub_991_2_n_114);
 assign sub_991_2_n_140 = ~(sub_991_2_n_132 & (sub_991_2_n_133 | sub_991_2_n_122));
 assign sub_991_2_n_139 = ~(sub_991_2_n_136 & sub_991_2_n_103);
 assign sub_991_2_n_138 = ~(sub_991_2_n_137 | sub_991_2_n_131);
 assign sub_991_2_n_137 = ~(sub_991_2_n_130 | sub_991_2_n_123);
 assign sub_991_2_n_136 = ~(sub_991_2_n_135 & sub_991_2_n_49);
 assign sub_991_2_n_135 = ~(sub_991_2_n_128 | (sub_991_2_n_69 & in1_113_0_));
 assign in1_115_1_ = ~(in1_113_0_ ^ (n_1587 ^ sub_991_2_n_69));
 assign sub_991_2_n_133 = ~(sub_991_2_n_127 | sub_991_2_n_119);
 assign sub_991_2_n_132 = ~(sub_991_2_n_121 | (sub_991_2_n_116 & sub_991_2_n_100));
 assign sub_991_2_n_131 = ~(sub_991_2_n_113 & ~(sub_991_2_n_118 & sub_991_2_n_109));
 assign sub_991_2_n_130 = ~(sub_991_2_n_112 | ~(sub_991_2_n_115 | sub_991_2_n_20));
 assign sub_991_2_n_129 = ~(sub_991_2_n_126 | sub_991_2_n_111);
 assign sub_991_2_n_128 = ~(n_1587 | ~sub_991_2_n_69);
 assign sub_991_2_n_127 = ~(sub_991_2_n_124 | sub_991_2_n_108);
 assign sub_991_2_n_126 = ~(sub_991_2_n_117 | sub_991_2_n_10);
 assign sub_991_2_n_125 = ~(sub_991_2_n_32 | sub_991_2_n_123);
 assign sub_991_2_n_121 = ~(sub_991_2_n_66 & (sub_991_2_n_57 | sub_991_2_n_74));
 assign sub_991_2_n_120 = ~(sub_991_2_n_97 | sub_991_2_n_108);
 assign sub_991_2_n_119 = ~(sub_991_2_n_65 & (sub_991_2_n_85 | sub_991_2_n_83));
 assign sub_991_2_n_124 = ~(sub_991_2_n_88 | ~(sub_991_2_n_53 | sub_991_2_n_51));
 assign sub_991_2_n_123 = ~(sub_991_2_n_98 & sub_991_2_n_109);
 assign sub_991_2_n_122 = ~(sub_991_2_n_94 & sub_991_2_n_100);
 assign sub_991_2_n_114 = ~(sub_991_2_n_104 | sub_991_2_n_62);
 assign sub_991_2_n_113 = ~(sub_991_2_n_63 | ~(sub_991_2_n_56 | sub_991_2_n_76));
 assign sub_991_2_n_112 = ~(sub_991_2_n_61 & (sub_991_2_n_75 | sub_991_2_n_6));
 assign sub_991_2_n_111 = ~(sub_991_2_n_64 & (sub_991_2_n_60 | sub_991_2_n_4));
 assign sub_991_2_n_118 = ~(sub_991_2_n_90 & (sub_991_2_n_81 | sub_991_2_n_0));
 assign sub_991_2_n_117 = ~(sub_991_2_n_67 | ~(sub_991_2_n_87 | sub_991_2_n_71));
 assign sub_991_2_n_116 = ~(sub_991_2_n_89 & (sub_991_2_n_52 | sub_991_2_n_59));
 assign sub_991_2_n_115 = ~(sub_991_2_n_68 | ~(sub_991_2_n_55 | sub_991_2_n_58));
 assign sub_991_2_n_104 = ~(sub_991_2_n_77 | sub_991_2_n_79);
 assign sub_991_2_n_103 = ~(sub_991_2_n_72 | sub_991_2_n_79);
 assign sub_991_2_n_102 = ~(sub_991_2_n_84 | sub_991_2_n_87);
 assign sub_991_2_n_110 = ~(sub_991_2_n_62 | sub_991_2_n_79);
 assign sub_991_2_n_109 = ~(sub_991_2_n_5 | sub_991_2_n_76);
 assign sub_991_2_n_108 = ~(sub_991_2_n_1 & ~sub_991_2_n_83);
 assign sub_991_2_n_107 = ~(sub_991_2_n_63 | sub_991_2_n_76);
 assign sub_991_2_n_106 = ~(sub_991_2_n_78 | sub_991_2_n_72);
 assign sub_991_2_n_105 = ~(sub_991_2_n_88 | sub_991_2_n_51);
 assign sub_991_2_n_96 = ~sub_991_2_n_95;
 assign in1_115_0_ = ~(sub_991_2_n_69 & ~(sub_991_2_n_48 & n_1510));
 assign sub_991_2_n_101 = ~(sub_991_2_n_6 | ~sub_991_2_n_61);
 assign sub_991_2_n_100 = ~(sub_991_2_n_2 | sub_991_2_n_74);
 assign sub_991_2_n_99 = ~(sub_991_2_n_68 | sub_991_2_n_58);
 assign sub_991_2_n_98 = ~(sub_991_2_n_3 | sub_991_2_n_0);
 assign sub_991_2_n_91 = (sub_991_2_n_67 | sub_991_2_n_87);
 assign sub_991_2_n_97 = (sub_991_2_n_70 | sub_991_2_n_51);
 assign sub_991_2_n_95 = ~(sub_991_2_n_82 | sub_991_2_n_58);
 assign sub_991_2_n_94 = ~(sub_991_2_n_50 | sub_991_2_n_59);
 assign sub_991_2_n_93 = ~(sub_991_2_n_74 | ~sub_991_2_n_66);
 assign sub_991_2_n_86 = ~sub_991_2_n_85;
 assign sub_991_2_n_78 = ~sub_991_2_n_77;
 assign sub_991_2_n_73 = ~sub_991_2_n_72;
 assign sub_991_2_n_90 = ~(in1_113_20_ & ~n_1594);
 assign sub_991_2_n_89 = ~(in1_113_12_ & ~n_1582);
 assign sub_991_2_n_88 = ~(n_1590 | ~in1_113_8_);
 assign sub_991_2_n_87 = ~(in1_113_4_ | ~n_1570);
 assign sub_991_2_n_85 = ~(in1_113_9_ & ~n_1552);
 assign sub_991_2_n_84 = ~(in1_113_3_ | ~n_1536);
 assign sub_991_2_n_83 = ~(in1_113_10_ | ~n_1556);
 assign sub_991_2_n_82 = ~(in1_113_15_ | ~n_1550);
 assign sub_991_2_n_81 = ~(in1_113_19_ & ~n_1566);
 assign sub_991_2_n_80 = ~(in1_113_5_ | ~n_1568);
 assign sub_991_2_n_79 = ~(in1_113_2_ | sub_991_2_n_47);
 assign sub_991_2_n_77 = ~(in1_113_1_ & ~n_1478);
 assign sub_991_2_n_76 = ~(in1_113_22_ | ~n_1404);
 assign sub_991_2_n_75 = ~(in1_113_17_ & ~n_1473);
 assign sub_991_2_n_74 = ~(in1_113_14_ | ~n_1496);
 assign sub_991_2_n_72 = ~(in1_113_1_ | ~n_1478);
 assign sub_991_2_n_71 = ~(in1_113_3_ & ~n_1536);
 assign sub_991_2_n_70 = ~(in1_113_7_ | ~n_1480);
 assign sub_991_2_n_69 = ~(n_1544 & ~n_1510);
 assign sub_991_2_n_49 = ~(in1_113_0_ & ~n_1587);
 assign sub_991_2_n_68 = ~(n_1563 | ~in1_113_16_);
 assign sub_991_2_n_67 = ~(n_1570 | ~in1_113_4_);
 assign sub_991_2_n_66 = ~(in1_113_14_ & ~n_1496);
 assign sub_991_2_n_65 = ~(in1_113_10_ & ~n_1556);
 assign sub_991_2_n_64 = ~(in1_113_6_ & ~n_1528);
 assign sub_991_2_n_63 = ~(n_1404 | ~in1_113_22_);
 assign sub_991_2_n_62 = (sub_991_2_n_47 & in1_113_2_);
 assign sub_991_2_n_61 = ~(in1_113_18_ & ~n_1559);
 assign sub_991_2_n_60 = ~(in1_113_5_ & ~n_1568);
 assign sub_991_2_n_59 = ~(in1_113_12_ | ~n_1582);
 assign sub_991_2_n_58 = ~(in1_113_16_ | ~n_1563);
 assign sub_991_2_n_57 = ~(in1_113_13_ & ~n_1578);
 assign sub_991_2_n_56 = ~(in1_113_21_ & ~n_1592);
 assign sub_991_2_n_55 = ~(in1_113_15_ & ~n_1550);
 assign sub_991_2_n_54 = ~(in1_113_17_ | ~n_1473);
 assign sub_991_2_n_53 = ~(in1_113_7_ & ~n_1480);
 assign sub_991_2_n_52 = ~(in1_113_11_ & ~n_1596);
 assign sub_991_2_n_51 = ~(in1_113_8_ | ~n_1590);
 assign sub_991_2_n_50 = ~(in1_113_11_ | ~n_1596);
 assign sub_991_2_n_48 = ~n_1544;
 assign sub_991_2_n_47 = ~n_1580;
 assign in1_115_14_ = ~(sub_991_2_n_159 ^ sub_991_2_n_12);
 assign in1_115_12_ = ~(sub_991_2_n_44 ^ sub_991_2_n_7);
 assign sub_991_2_n_44 = (sub_991_2_n_151 & sub_991_2_n_133);
 assign sub_991_2_n_43 = (sub_991_2_n_145 & sub_991_2_n_117);
 assign in1_115_20_ = (sub_991_2_n_166 ^ sub_991_2_n_19);
 assign in1_115_10_ = (sub_991_2_n_153 ^ sub_991_2_n_17);
 assign in1_115_3_ = ~(sub_991_2_n_143 ^ sub_991_2_n_110);
 assign in1_115_7_ = (sub_991_2_n_150 ^ sub_991_2_n_14);
 assign in1_115_23_ = (sub_991_2_n_172 ^ sub_991_2_n_107);
 assign in1_115_2_ = (sub_991_2_n_136 ^ sub_991_2_n_106);
 assign in1_115_4_ = ~(sub_991_2_n_142 ^ sub_991_2_n_16);
 assign in1_115_22_ = ~(sub_991_2_n_171 ^ sub_991_2_n_11);
 assign in1_115_21_ = (sub_991_2_n_170 ^ sub_991_2_n_22);
 assign in1_115_9_ = (sub_991_2_n_152 ^ sub_991_2_n_105);
 assign sub_991_2_n_32 = ~(sub_991_2_n_95 & ~sub_991_2_n_20);
 assign in1_115_19_ = (sub_991_2_n_169 ^ sub_991_2_n_101);
 assign in1_115_8_ = (sub_991_2_n_148 ^ sub_991_2_n_8);
 assign in1_115_18_ = (sub_991_2_n_163 ^ sub_991_2_n_18);
 assign in1_115_17_ = (sub_991_2_n_162 ^ sub_991_2_n_99);
 assign in1_115_6_ = ~(sub_991_2_n_43 ^ sub_991_2_n_13);
 assign in1_115_13_ = (sub_991_2_n_158 ^ sub_991_2_n_21);
 assign sub_991_2_n_25 = ~(sub_991_2_n_44 | ~sub_991_2_n_94);
 assign in1_115_11_ = ~(sub_991_2_n_157 ^ sub_991_2_n_15);
 assign in1_115_15_ = (sub_991_2_n_167 ^ sub_991_2_n_93);
 assign sub_991_2_n_22 = ~(sub_991_2_n_0 | ~sub_991_2_n_90);
 assign sub_991_2_n_21 = ~(sub_991_2_n_59 | ~sub_991_2_n_89);
 assign sub_991_2_n_20 = (sub_991_2_n_6 | sub_991_2_n_54);
 assign sub_991_2_n_19 = ~(sub_991_2_n_3 | ~sub_991_2_n_81);
 assign sub_991_2_n_18 = ~(sub_991_2_n_54 | ~sub_991_2_n_75);
 assign sub_991_2_n_17 = ~(sub_991_2_n_86 | ~sub_991_2_n_1);
 assign sub_991_2_n_16 = ~(sub_991_2_n_84 | ~sub_991_2_n_71);
 assign sub_991_2_n_15 = ~(sub_991_2_n_83 | ~sub_991_2_n_65);
 assign sub_991_2_n_14 = ~(sub_991_2_n_4 | ~sub_991_2_n_64);
 assign sub_991_2_n_13 = ~(sub_991_2_n_80 | ~sub_991_2_n_60);
 assign sub_991_2_n_12 = ~(sub_991_2_n_2 | ~sub_991_2_n_57);
 assign sub_991_2_n_11 = ~(sub_991_2_n_5 | ~sub_991_2_n_56);
 assign sub_991_2_n_10 = (sub_991_2_n_4 | sub_991_2_n_80);
 assign sub_991_2_n_9 = ~(sub_991_2_n_82 | ~sub_991_2_n_55);
 assign sub_991_2_n_8 = ~(sub_991_2_n_70 | ~sub_991_2_n_53);
 assign sub_991_2_n_7 = ~(sub_991_2_n_50 | ~sub_991_2_n_52);
 assign sub_991_2_n_6 = ~(in1_113_18_ | ~n_1559);
 assign sub_991_2_n_5 = ~(in1_113_21_ | ~n_1592);
 assign sub_991_2_n_4 = ~(in1_113_6_ | ~n_1528);
 assign sub_991_2_n_3 = ~(in1_113_19_ | ~n_1566);
 assign sub_991_2_n_2 = ~(in1_113_13_ | ~n_1578);
 assign sub_991_2_n_1 = ~(n_1552 & ~in1_113_9_);
 assign sub_991_2_n_0 = ~(in1_113_20_ | ~n_1594);
 assign sub_1012_2_n_188 = ~(sub_1012_2_n_50 | ~(sub_1012_2_n_187 | sub_1012_2_n_51));
 assign sub_1012_2_n_186 = ~(sub_1012_2_n_180 | sub_1012_2_n_75);
 assign sub_1012_2_n_185 = ~(sub_1012_2_n_179 | sub_1012_2_n_39);
 assign sub_1012_2_n_184 = ~(sub_1012_2_n_178 | sub_1012_2_n_41);
 assign sub_1012_2_n_187 = ~(sub_1012_2_n_181 | sub_1012_2_n_118);
 assign in1_118_14_ = ~(sub_1012_2_n_24 ^ sub_1012_2_n_90);
 assign in1_118_13_ = ~(sub_1012_2_n_170 ^ sub_1012_2_n_88);
 assign sub_1012_2_n_181 = ~(sub_1012_2_n_176 | sub_1012_2_n_94);
 assign sub_1012_2_n_180 = ~(sub_1012_2_n_176 | sub_1012_2_n_69);
 assign sub_1012_2_n_179 = ~(sub_1012_2_n_177 | sub_1012_2_n_38);
 assign sub_1012_2_n_178 = ~(sub_1012_2_n_24 | sub_1012_2_n_46);
 assign sub_1012_2_n_175 = ~(sub_1012_2_n_163 & sub_1012_2_n_148);
 assign sub_1012_2_n_174 = ~(sub_1012_2_n_167 | sub_1012_2_n_37);
 assign sub_1012_2_n_177 = ~(sub_1012_2_n_23 | sub_1012_2_n_119);
 assign sub_1012_2_n_176 = ~(sub_1012_2_n_168 | sub_1012_2_n_136);
 assign in1_118_10_ = ~(sub_1012_2_n_160 ^ sub_1012_2_n_86);
 assign in1_118_12_ = ~(sub_1012_2_n_161 ^ sub_1012_2_n_89);
 assign in1_118_9_ = ~(sub_1012_2_n_159 ^ sub_1012_2_n_8);
 assign sub_1012_2_n_170 = ~(sub_1012_2_n_165 | sub_1012_2_n_45);
 assign sub_1012_2_n_169 = ~(sub_1012_2_n_164 | sub_1012_2_n_63);
 assign sub_1012_2_n_168 = ~(sub_1012_2_n_162 | sub_1012_2_n_124);
 assign sub_1012_2_n_167 = ~(sub_1012_2_n_162 | sub_1012_2_n_72);
 assign sub_1012_2_n_166 = ~(sub_1012_2_n_161 | sub_1012_2_n_7);
 assign sub_1012_2_n_165 = ~(sub_1012_2_n_161 | sub_1012_2_n_60);
 assign sub_1012_2_n_164 = ~(sub_1012_2_n_160 | sub_1012_2_n_66);
 assign sub_1012_2_n_163 = ~(sub_1012_2_n_142 | (sub_1012_2_n_156 & sub_1012_2_n_25));
 assign sub_1012_2_n_162 = ~(sub_1012_2_n_156 | sub_1012_2_n_144);
 assign sub_1012_2_n_161 = ~(sub_1012_2_n_135 | ~(sub_1012_2_n_154 | sub_1012_2_n_126));
 assign sub_1012_2_n_160 = ~(sub_1012_2_n_157 | sub_1012_2_n_127);
 assign sub_1012_2_n_159 = ~(sub_1012_2_n_79 | ~(sub_1012_2_n_154 | sub_1012_2_n_43));
 assign in1_118_8_ = ~(sub_1012_2_n_154 ^ sub_1012_2_n_87);
 assign sub_1012_2_n_157 = ~(sub_1012_2_n_154 | sub_1012_2_n_93);
 assign sub_1012_2_n_156 = ~(sub_1012_2_n_154 | sub_1012_2_n_131);
 assign sub_1012_2_n_155 = ~(sub_1012_2_n_62 | (sub_1012_2_n_152 & sub_1012_2_n_0));
 assign sub_1012_2_n_154 = ~(sub_1012_2_n_153 | sub_1012_2_n_134);
 assign sub_1012_2_n_153 = ~(sub_1012_2_n_149 | sub_1012_2_n_95);
 assign sub_1012_2_n_152 = ~(sub_1012_2_n_149 & sub_1012_2_n_121);
 assign sub_1012_2_n_151 = ~(sub_1012_2_n_31 | (sub_1012_2_n_145 & sub_1012_2_n_34));
 assign in1_118_4_ = (sub_1012_2_n_145 ^ sub_1012_2_n_91);
 assign sub_1012_2_n_149 = ~(sub_1012_2_n_145 & sub_1012_2_n_101);
 assign sub_1012_2_n_148 = ~(sub_1012_2_n_144 & sub_1012_2_n_25);
 assign sub_1012_2_n_147 = ~(sub_1012_2_n_48 | (sub_1012_2_n_141 & sub_1012_2_n_65));
 assign in1_118_2_ = (sub_1012_2_n_141 ^ sub_1012_2_n_100);
 assign sub_1012_2_n_145 = ~(sub_1012_2_n_143 & sub_1012_2_n_123);
 assign sub_1012_2_n_144 = ~(sub_1012_2_n_138 & ~(sub_1012_2_n_135 & sub_1012_2_n_129));
 assign sub_1012_2_n_143 = ~(sub_1012_2_n_141 & sub_1012_2_n_102);
 assign sub_1012_2_n_142 = ~(sub_1012_2_n_137 & ~(sub_1012_2_n_136 & sub_1012_2_n_128));
 assign sub_1012_2_n_141 = ~(sub_1012_2_n_140 & sub_1012_2_n_56);
 assign sub_1012_2_n_140 = ~(sub_1012_2_n_133 | (sub_1012_2_n_130 & in1_116_0_));
 assign in1_118_1_ = ~((sub_1012_2_n_58 & ~sub_1012_2_n_5) | (sub_1012_2_n_130 & sub_1012_2_n_5));
 assign sub_1012_2_n_138 = ~(sub_1012_2_n_132 | sub_1012_2_n_114);
 assign sub_1012_2_n_137 = ~(sub_1012_2_n_116 | (sub_1012_2_n_118 & sub_1012_2_n_109));
 assign sub_1012_2_n_136 = ~(sub_1012_2_n_117 & ~(sub_1012_2_n_119 & sub_1012_2_n_105));
 assign sub_1012_2_n_135 = ~(sub_1012_2_n_122 & ~(sub_1012_2_n_127 & sub_1012_2_n_110));
 assign sub_1012_2_n_134 = ~(sub_1012_2_n_115 & (sub_1012_2_n_121 | sub_1012_2_n_95));
 assign sub_1012_2_n_133 = ~(sub_1012_2_n_58 | n_1587);
 assign sub_1012_2_n_132 = ~(sub_1012_2_n_120 | sub_1012_2_n_99);
 assign sub_1012_2_n_131 = ~(sub_1012_2_n_125 & sub_1012_2_n_129);
 assign sub_1012_2_n_130 = ~sub_1012_2_n_58;
 assign sub_1012_2_n_126 = ~sub_1012_2_n_125;
 assign sub_1012_2_n_123 = ~(sub_1012_2_n_81 | ~(sub_1012_2_n_47 | sub_1012_2_n_68));
 assign sub_1012_2_n_122 = ~(sub_1012_2_n_84 | (sub_1012_2_n_63 & sub_1012_2_n_32));
 assign sub_1012_2_n_129 = ~(sub_1012_2_n_7 | sub_1012_2_n_99);
 assign sub_1012_2_n_128 = ~(sub_1012_2_n_94 | ~sub_1012_2_n_109);
 assign sub_1012_2_n_127 = ~(sub_1012_2_n_80 & (sub_1012_2_n_78 | sub_1012_2_n_59));
 assign sub_1012_2_n_125 = ~(sub_1012_2_n_93 | ~sub_1012_2_n_110);
 assign sub_1012_2_n_124 = ~(sub_1012_2_n_113 & sub_1012_2_n_105);
 assign sub_1012_2_n_117 = ~(sub_1012_2_n_57 | (sub_1012_2_n_39 & sub_1012_2_n_76));
 assign sub_1012_2_n_116 = ~(sub_1012_2_n_53 & (sub_1012_2_n_49 | sub_1012_2_n_67));
 assign sub_1012_2_n_115 = ~(sub_1012_2_n_82 | ~(sub_1012_2_n_61 | sub_1012_2_n_35));
 assign sub_1012_2_n_114 = ~(sub_1012_2_n_54 & ~(sub_1012_2_n_41 & sub_1012_2_n_71));
 assign sub_1012_2_n_121 = ~(sub_1012_2_n_55 | ~(sub_1012_2_n_30 | sub_1012_2_n_70));
 assign sub_1012_2_n_120 = ~(sub_1012_2_n_85 | ~(sub_1012_2_n_44 | sub_1012_2_n_73));
 assign sub_1012_2_n_119 = ~(sub_1012_2_n_52 & (sub_1012_2_n_36 | sub_1012_2_n_42));
 assign sub_1012_2_n_118 = ~(sub_1012_2_n_83 & (sub_1012_2_n_74 | sub_1012_2_n_40));
 assign sub_1012_2_n_102 = ~(sub_1012_2_n_64 | sub_1012_2_n_68);
 assign sub_1012_2_n_101 = ~(sub_1012_2_n_33 | sub_1012_2_n_70);
 assign sub_1012_2_n_113 = ~(sub_1012_2_n_72 | sub_1012_2_n_42);
 assign sub_1012_2_n_112 = ~(sub_1012_2_n_81 | sub_1012_2_n_68);
 assign sub_1012_2_n_111 = ~(sub_1012_2_n_55 | sub_1012_2_n_70);
 assign sub_1012_2_n_100 = ~(sub_1012_2_n_48 | sub_1012_2_n_64);
 assign sub_1012_2_n_110 = ~(sub_1012_2_n_66 | sub_1012_2_n_2);
 assign sub_1012_2_n_109 = ~(sub_1012_2_n_51 | sub_1012_2_n_67);
 assign sub_1012_2_n_108 = ~(sub_1012_2_n_53 & ~sub_1012_2_n_67);
 assign sub_1012_2_n_107 = ~(sub_1012_2_n_50 | sub_1012_2_n_51);
 assign sub_1012_2_n_106 = ~(sub_1012_2_n_82 | sub_1012_2_n_35);
 assign sub_1012_2_n_105 = ~(sub_1012_2_n_38 | sub_1012_2_n_77);
 assign sub_1012_2_n_104 = ~(sub_1012_2_n_75 | sub_1012_2_n_69);
 assign sub_1012_2_n_103 = ~(sub_1012_2_n_57 | sub_1012_2_n_77);
 assign in1_118_0_ = ~(sub_1012_2_n_130 & ~(sub_1012_2_n_28 & n_1547));
 assign sub_1012_2_n_99 = ~(sub_1012_2_n_71 & ~sub_1012_2_n_46);
 assign sub_1012_2_n_98 = ~(sub_1012_2_n_39 | sub_1012_2_n_38);
 assign sub_1012_2_n_91 = ~(sub_1012_2_n_31 | sub_1012_2_n_33);
 assign sub_1012_2_n_97 = ~(sub_1012_2_n_37 | sub_1012_2_n_72);
 assign sub_1012_2_n_96 = ~(sub_1012_2_n_84 | sub_1012_2_n_2);
 assign sub_1012_2_n_90 = ~(sub_1012_2_n_41 | sub_1012_2_n_46);
 assign sub_1012_2_n_89 = ~(sub_1012_2_n_45 | sub_1012_2_n_60);
 assign sub_1012_2_n_88 = ~(sub_1012_2_n_85 | sub_1012_2_n_73);
 assign sub_1012_2_n_95 = ~(sub_1012_2_n_0 & ~sub_1012_2_n_35);
 assign sub_1012_2_n_87 = ~(sub_1012_2_n_79 | sub_1012_2_n_43);
 assign sub_1012_2_n_86 = ~(sub_1012_2_n_63 | sub_1012_2_n_66);
 assign sub_1012_2_n_94 = (sub_1012_2_n_69 | sub_1012_2_n_40);
 assign sub_1012_2_n_93 = (sub_1012_2_n_43 | sub_1012_2_n_59);
 assign sub_1012_2_n_79 = ~sub_1012_2_n_78;
 assign sub_1012_2_n_76 = ~sub_1012_2_n_77;
 assign sub_1012_2_n_75 = ~sub_1012_2_n_74;
 assign sub_1012_2_n_65 = ~sub_1012_2_n_64;
 assign sub_1012_2_n_62 = ~sub_1012_2_n_61;
 assign sub_1012_2_n_85 = ~(n_1582 | ~in1_116_12_);
 assign sub_1012_2_n_84 = ~(n_1556 | ~in1_116_10_);
 assign sub_1012_2_n_83 = ~(in1_116_20_ & ~n_1594);
 assign sub_1012_2_n_82 = ~(n_1528 | ~in1_116_6_);
 assign sub_1012_2_n_81 = ~(n_1580 | ~in1_116_2_);
 assign sub_1012_2_n_80 = ~(in1_116_8_ & ~n_1590);
 assign sub_1012_2_n_78 = ~(in1_116_7_ & ~n_1480);
 assign sub_1012_2_n_77 = ~(in1_116_18_ | sub_1012_2_n_27);
 assign sub_1012_2_n_74 = ~(in1_116_19_ & ~n_1566);
 assign sub_1012_2_n_73 = ~(in1_116_12_ | ~n_1582);
 assign sub_1012_2_n_72 = ~(in1_116_15_ | ~n_1550);
 assign sub_1012_2_n_71 = ~(n_1496 & ~in1_116_14_);
 assign sub_1012_2_n_70 = ~(in1_116_4_ | ~n_1570);
 assign sub_1012_2_n_69 = ~(in1_116_19_ | ~n_1566);
 assign sub_1012_2_n_68 = ~(in1_116_2_ | ~n_1580);
 assign sub_1012_2_n_67 = ~(in1_116_22_ | ~n_1404);
 assign sub_1012_2_n_66 = ~(in1_116_9_ | ~n_1552);
 assign sub_1012_2_n_64 = ~(in1_116_1_ | ~n_1478);
 assign sub_1012_2_n_63 = ~(n_1552 | ~in1_116_9_);
 assign sub_1012_2_n_61 = ~(in1_116_5_ & ~n_1568);
 assign sub_1012_2_n_60 = ~(in1_116_11_ | ~n_1596);
 assign sub_1012_2_n_59 = ~(in1_116_8_ | ~n_1590);
 assign sub_1012_2_n_58 = ~(n_1547 | sub_1012_2_n_28);
 assign sub_1012_2_n_50 = ~sub_1012_2_n_49;
 assign sub_1012_2_n_48 = ~sub_1012_2_n_47;
 assign sub_1012_2_n_45 = ~sub_1012_2_n_44;
 assign sub_1012_2_n_37 = ~sub_1012_2_n_36;
 assign sub_1012_2_n_34 = ~sub_1012_2_n_33;
 assign sub_1012_2_n_32 = ~sub_1012_2_n_2;
 assign sub_1012_2_n_31 = ~sub_1012_2_n_30;
 assign sub_1012_2_n_29 = ~(in1_116_0_ | ~n_1587);
 assign sub_1012_2_n_57 = (sub_1012_2_n_27 & in1_116_18_);
 assign sub_1012_2_n_56 = ~(in1_116_0_ & ~n_1587);
 assign sub_1012_2_n_55 = ~(n_1570 | ~in1_116_4_);
 assign sub_1012_2_n_54 = ~(in1_116_14_ & ~n_1496);
 assign sub_1012_2_n_53 = ~(in1_116_22_ & ~n_1404);
 assign sub_1012_2_n_52 = ~(in1_116_16_ & ~n_1563);
 assign sub_1012_2_n_51 = ~(in1_116_21_ | ~n_1592);
 assign sub_1012_2_n_49 = ~(in1_116_21_ & ~n_1592);
 assign sub_1012_2_n_47 = ~(in1_116_1_ & ~n_1478);
 assign sub_1012_2_n_46 = ~(in1_116_13_ | ~n_1578);
 assign sub_1012_2_n_44 = ~(in1_116_11_ & ~n_1596);
 assign sub_1012_2_n_43 = ~(in1_116_7_ | ~n_1480);
 assign sub_1012_2_n_42 = ~(in1_116_16_ | ~n_1563);
 assign sub_1012_2_n_41 = ~(n_1578 | ~in1_116_13_);
 assign sub_1012_2_n_40 = ~(in1_116_20_ | ~n_1594);
 assign sub_1012_2_n_39 = ~(n_1473 | ~in1_116_17_);
 assign sub_1012_2_n_38 = ~(in1_116_17_ | ~n_1473);
 assign sub_1012_2_n_36 = ~(in1_116_15_ & ~n_1550);
 assign sub_1012_2_n_35 = ~(in1_116_6_ | ~n_1528);
 assign sub_1012_2_n_33 = ~(in1_116_3_ | ~n_1536);
 assign sub_1012_2_n_30 = ~(in1_116_3_ & ~n_1536);
 assign sub_1012_2_n_28 = ~n_1544;
 assign sub_1012_2_n_27 = ~n_1559;
 assign in1_118_6_ = (sub_1012_2_n_152 ^ sub_1012_2_n_3);
 assign sub_1012_2_n_25 = ~(sub_1012_2_n_124 | ~sub_1012_2_n_128);
 assign sub_1012_2_n_24 = ~(sub_1012_2_n_166 | ~sub_1012_2_n_120);
 assign sub_1012_2_n_23 = ~(sub_1012_2_n_162 | ~sub_1012_2_n_113);
 assign in1_118_3_ = ~(sub_1012_2_n_147 ^ sub_1012_2_n_112);
 assign in1_118_5_ = ~(sub_1012_2_n_151 ^ sub_1012_2_n_111);
 assign in1_118_23_ = (sub_1012_2_n_188 ^ sub_1012_2_n_108);
 assign in1_118_22_ = ~(sub_1012_2_n_187 ^ sub_1012_2_n_107);
 assign in1_118_21_ = ~(sub_1012_2_n_186 ^ sub_1012_2_n_9);
 assign in1_118_7_ = ~(sub_1012_2_n_155 ^ sub_1012_2_n_106);
 assign in1_118_20_ = ~(sub_1012_2_n_176 ^ sub_1012_2_n_104);
 assign in1_118_19_ = ~(sub_1012_2_n_185 ^ sub_1012_2_n_103);
 assign in1_118_18_ = ~(sub_1012_2_n_177 ^ sub_1012_2_n_98);
 assign in1_118_17_ = ~(sub_1012_2_n_174 ^ sub_1012_2_n_4);
 assign in1_118_16_ = ~(sub_1012_2_n_162 ^ sub_1012_2_n_97);
 assign in1_118_11_ = ~(sub_1012_2_n_169 ^ sub_1012_2_n_96);
 assign in1_118_15_ = ~(sub_1012_2_n_184 ^ sub_1012_2_n_6);
 assign sub_1012_2_n_9 = ~(sub_1012_2_n_40 | ~sub_1012_2_n_83);
 assign sub_1012_2_n_8 = ~(sub_1012_2_n_59 | ~sub_1012_2_n_80);
 assign sub_1012_2_n_7 = (sub_1012_2_n_73 | sub_1012_2_n_60);
 assign sub_1012_2_n_6 = (sub_1012_2_n_54 & sub_1012_2_n_71);
 assign sub_1012_2_n_5 = ~(sub_1012_2_n_29 | ~sub_1012_2_n_56);
 assign sub_1012_2_n_4 = ~(sub_1012_2_n_42 | ~sub_1012_2_n_52);
 assign sub_1012_2_n_3 = ~(sub_1012_2_n_62 | ~sub_1012_2_n_0);
 assign sub_1012_2_n_2 = ~(in1_116_10_ | ~n_1556);
 assign in1_118_24_ = ~(sub_1012_2_n_175 ^ in1_116_23_);
 assign sub_1012_2_n_0 = ~(n_1568 & ~in1_116_5_);
 assign sub_1033_2_n_167 = ~(sub_1033_2_n_43 & (sub_1033_2_n_166 | sub_1033_2_n_40));
 assign sub_1033_2_n_166 = ~sub_1033_2_n_165;
 assign sub_1033_2_n_165 = ~(sub_1033_2_n_106 & (sub_1033_2_n_158 | sub_1033_2_n_83));
 assign sub_1033_2_n_164 = ~(sub_1033_2_n_65 & (sub_1033_2_n_158 | sub_1033_2_n_64));
 assign sub_1033_2_n_163 = ~(sub_1033_2_n_71 & (sub_1033_2_n_157 | sub_1033_2_n_45));
 assign in1_121_20_ = (sub_1033_2_n_158 ^ sub_1033_2_n_89);
 assign in1_121_18_ = (sub_1033_2_n_157 ^ sub_1033_2_n_88);
 assign sub_1033_2_n_160 = ~(sub_1033_2_n_39 & (sub_1033_2_n_152 | sub_1033_2_n_50));
 assign in1_121_24_ = ~(sub_1033_2_n_153 ^ in1_119_23_);
 assign sub_1033_2_n_158 = ~(sub_1033_2_n_154 | sub_1033_2_n_121);
 assign sub_1033_2_n_157 = ~(sub_1033_2_n_16 | sub_1033_2_n_107);
 assign sub_1033_2_n_156 = ~(sub_1033_2_n_69 & (sub_1033_2_n_32 | sub_1033_2_n_42));
 assign in1_121_16_ = (sub_1033_2_n_32 ^ sub_1033_2_n_79);
 assign sub_1033_2_n_154 = ~(sub_1033_2_n_32 | sub_1033_2_n_110);
 assign sub_1033_2_n_153 = ~(sub_1033_2_n_134 & (sub_1033_2_n_147 | sub_1033_2_n_114));
 assign sub_1033_2_n_152 = ~(sub_1033_2_n_149 | sub_1033_2_n_111);
 assign sub_1033_2_n_151 = ~(sub_1033_2_n_70 & (sub_1033_2_n_146 | sub_1033_2_n_46));
 assign in1_121_12_ = ~(sub_1033_2_n_146 ^ sub_1033_2_n_10);
 assign sub_1033_2_n_149 = ~(sub_1033_2_n_146 | sub_1033_2_n_93);
 assign sub_1033_2_n_148 = ~(sub_1033_2_n_61 & (sub_1033_2_n_31 | sub_1033_2_n_1));
 assign sub_1033_2_n_147 = ~(sub_1033_2_n_22 & sub_1033_2_n_29);
 assign sub_1033_2_n_146 = ~(sub_1033_2_n_22 | sub_1033_2_n_119);
 assign sub_1033_2_n_145 = ~(sub_1033_2_n_48 & (sub_1033_2_n_140 | sub_1033_2_n_47));
 assign in1_121_8_ = ~(sub_1033_2_n_140 ^ sub_1033_2_n_4);
 assign sub_1033_2_n_143 = ~(sub_1033_2_n_63 & (sub_1033_2_n_138 | sub_1033_2_n_68));
 assign sub_1033_2_n_142 = ~(sub_1033_2_n_139 & sub_1033_2_n_81);
 assign in1_121_5_ = (sub_1033_2_n_136 ^ sub_1033_2_n_7);
 assign sub_1033_2_n_140 = ~sub_1033_2_n_139;
 assign sub_1033_2_n_139 = ~(sub_1033_2_n_137 & sub_1033_2_n_120);
 assign sub_1033_2_n_138 = ~(sub_1033_2_n_135 | sub_1033_2_n_105);
 assign sub_1033_2_n_137 = ~(sub_1033_2_n_135 & sub_1033_2_n_97);
 assign sub_1033_2_n_136 = ~(sub_1033_2_n_73 & (sub_1033_2_n_130 | sub_1033_2_n_59));
 assign sub_1033_2_n_135 = ~(sub_1033_2_n_130 | sub_1033_2_n_90);
 assign sub_1033_2_n_134 = ~(sub_1033_2_n_133 | sub_1033_2_n_125);
 assign sub_1033_2_n_133 = ~(sub_1033_2_n_126 | sub_1033_2_n_114);
 assign sub_1033_2_n_132 = ~(sub_1033_2_n_44 & (sub_1033_2_n_123 | sub_1033_2_n_66));
 assign in1_121_2_ = ~(sub_1033_2_n_129 & ~sub_1033_2_n_128);
 assign sub_1033_2_n_130 = ~(sub_1033_2_n_127 | sub_1033_2_n_102);
 assign sub_1033_2_n_129 = ~(sub_1033_2_n_124 & sub_1033_2_n_100);
 assign sub_1033_2_n_128 = ~(sub_1033_2_n_124 | sub_1033_2_n_100);
 assign sub_1033_2_n_127 = ~(sub_1033_2_n_123 | sub_1033_2_n_11);
 assign sub_1033_2_n_126 = ~(sub_1033_2_n_118 | (sub_1033_2_n_119 & sub_1033_2_n_29));
 assign sub_1033_2_n_125 = ~(sub_1033_2_n_117 & ~(sub_1033_2_n_121 & sub_1033_2_n_113));
 assign sub_1033_2_n_123 = ~sub_1033_2_n_124;
 assign sub_1033_2_n_124 = ((sub_1033_2_n_36 & in1_119_0_) | ((in1_119_0_ & sub_1033_2_n_34) | (sub_1033_2_n_34
    & sub_1033_2_n_36)));
 assign in1_121_1_ = (in1_119_0_ ^ (sub_1033_2_n_34 ^ sub_1033_2_n_36));
 assign sub_1033_2_n_121 = ~(sub_1033_2_n_103 & ~(sub_1033_2_n_107 & sub_1033_2_n_92));
 assign sub_1033_2_n_120 = ~(sub_1033_2_n_104 | (sub_1033_2_n_105 & sub_1033_2_n_97));
 assign sub_1033_2_n_119 = ~(sub_1033_2_n_116 & sub_1033_2_n_108);
 assign sub_1033_2_n_118 = ~(sub_1033_2_n_109 & ~(sub_1033_2_n_111 & sub_1033_2_n_98));
 assign sub_1033_2_n_117 = ~(sub_1033_2_n_115 | sub_1033_2_n_101);
 assign sub_1033_2_n_116 = ~(sub_1033_2_n_112 & sub_1033_2_n_87);
 assign sub_1033_2_n_115 = ~(sub_1033_2_n_106 | sub_1033_2_n_96);
 assign sub_1033_2_n_114 = ~(sub_1033_2_n_113 & ~sub_1033_2_n_110);
 assign sub_1033_2_n_109 = ~(sub_1033_2_n_56 | ~(sub_1033_2_n_39 | sub_1033_2_n_60));
 assign sub_1033_2_n_108 = ~(sub_1033_2_n_74 | ~(sub_1033_2_n_61 | sub_1033_2_n_51));
 assign sub_1033_2_n_113 = ~(sub_1033_2_n_83 | sub_1033_2_n_96);
 assign sub_1033_2_n_112 = ~(sub_1033_2_n_52 & (sub_1033_2_n_48 | sub_1033_2_n_0));
 assign sub_1033_2_n_111 = ~(sub_1033_2_n_54 & (sub_1033_2_n_70 | sub_1033_2_n_41));
 assign sub_1033_2_n_110 = ~(sub_1033_2_n_84 & sub_1033_2_n_92);
 assign sub_1033_2_n_104 = ~(sub_1033_2_n_75 & (sub_1033_2_n_63 | sub_1033_2_n_58));
 assign sub_1033_2_n_103 = ~(sub_1033_2_n_77 | ~(sub_1033_2_n_71 | sub_1033_2_n_49));
 assign sub_1033_2_n_102 = ~(sub_1033_2_n_78 & (sub_1033_2_n_44 | sub_1033_2_n_72));
 assign sub_1033_2_n_101 = ~(sub_1033_2_n_55 & (sub_1033_2_n_43 | sub_1033_2_n_67));
 assign sub_1033_2_n_107 = ~(sub_1033_2_n_76 & (sub_1033_2_n_69 | sub_1033_2_n_37));
 assign sub_1033_2_n_106 = ~(sub_1033_2_n_53 | ~(sub_1033_2_n_65 | sub_1033_2_n_62));
 assign sub_1033_2_n_105 = ~(sub_1033_2_n_57 & (sub_1033_2_n_73 | sub_1033_2_n_38));
 assign sub_1033_2_n_90 = (sub_1033_2_n_59 | sub_1033_2_n_38);
 assign sub_1033_2_n_100 = ~(sub_1033_2_n_44 & ~sub_1033_2_n_66);
 assign sub_1033_2_n_99 = ~(sub_1033_2_n_67 | ~sub_1033_2_n_55);
 assign sub_1033_2_n_98 = ~(sub_1033_2_n_50 | sub_1033_2_n_60);
 assign sub_1033_2_n_97 = ~(sub_1033_2_n_68 | sub_1033_2_n_58);
 assign sub_1033_2_n_96 = (sub_1033_2_n_40 | sub_1033_2_n_67);
 assign sub_1033_2_n_95 = ~(sub_1033_2_n_53 | sub_1033_2_n_62);
 assign sub_1033_2_n_94 = ~(sub_1033_2_n_74 | sub_1033_2_n_51);
 assign sub_1033_2_n_93 = (sub_1033_2_n_46 | sub_1033_2_n_41);
 assign sub_1033_2_n_92 = ~(sub_1033_2_n_45 | sub_1033_2_n_49);
 assign sub_1033_2_n_89 = ~(sub_1033_2_n_65 & ~sub_1033_2_n_64);
 assign sub_1033_2_n_91 = ~(sub_1033_2_n_77 | sub_1033_2_n_49);
 assign sub_1033_2_n_88 = ~(sub_1033_2_n_71 & ~sub_1033_2_n_45);
 assign sub_1033_2_n_81 = ~(sub_1033_2_n_47 | sub_1033_2_n_0);
 assign in1_121_0_ = ~(sub_1033_2_n_36 & ~(sub_1033_2_n_35 & n_1402));
 assign sub_1033_2_n_87 = ~(sub_1033_2_n_1 | sub_1033_2_n_51);
 assign sub_1033_2_n_86 = ~(sub_1033_2_n_58 | ~sub_1033_2_n_75);
 assign sub_1033_2_n_85 = ~(sub_1033_2_n_56 | sub_1033_2_n_60);
 assign sub_1033_2_n_79 = ~(sub_1033_2_n_69 & ~sub_1033_2_n_42);
 assign sub_1033_2_n_84 = ~(sub_1033_2_n_42 | sub_1033_2_n_37);
 assign sub_1033_2_n_83 = (sub_1033_2_n_64 | sub_1033_2_n_62);
 assign sub_1033_2_n_82 = ~(sub_1033_2_n_37 | ~sub_1033_2_n_76);
 assign sub_1033_2_n_78 = ~(in1_119_2_ & ~n_1580);
 assign sub_1033_2_n_77 = ~(n_1559 | ~in1_119_18_);
 assign sub_1033_2_n_76 = ~(in1_119_16_ & ~n_1563);
 assign sub_1033_2_n_75 = ~(in1_119_6_ & ~n_1528);
 assign sub_1033_2_n_74 = ~(n_1556 | ~in1_119_10_);
 assign sub_1033_2_n_73 = ~(in1_119_3_ & ~n_1536);
 assign sub_1033_2_n_72 = ~(in1_119_2_ | ~n_1580);
 assign sub_1033_2_n_71 = ~(in1_119_17_ & ~n_1473);
 assign sub_1033_2_n_70 = ~(in1_119_11_ & ~n_1596);
 assign sub_1033_2_n_69 = ~(in1_119_15_ & ~n_1550);
 assign sub_1033_2_n_68 = ~(in1_119_5_ | ~n_1568);
 assign sub_1033_2_n_67 = ~(in1_119_22_ | ~n_1404);
 assign sub_1033_2_n_66 = ~(in1_119_1_ | ~n_1478);
 assign sub_1033_2_n_65 = ~(in1_119_19_ & ~n_1566);
 assign sub_1033_2_n_64 = ~(in1_119_19_ | ~n_1566);
 assign sub_1033_2_n_63 = ~(in1_119_5_ & ~n_1568);
 assign sub_1033_2_n_62 = ~(in1_119_20_ | ~n_1594);
 assign sub_1033_2_n_61 = ~(in1_119_9_ & ~n_1552);
 assign sub_1033_2_n_60 = ~(in1_119_14_ | ~n_1496);
 assign sub_1033_2_n_59 = ~(in1_119_3_ | ~n_1536);
 assign sub_1033_2_n_58 = ~(in1_119_6_ | ~n_1528);
 assign sub_1033_2_n_57 = ~(in1_119_4_ & ~n_1570);
 assign sub_1033_2_n_56 = ~(n_1496 | ~in1_119_14_);
 assign sub_1033_2_n_55 = ~(in1_119_22_ & ~n_1404);
 assign sub_1033_2_n_54 = ~(in1_119_12_ & ~n_1582);
 assign sub_1033_2_n_53 = ~(n_1594 | ~in1_119_20_);
 assign sub_1033_2_n_52 = ~(in1_119_8_ & ~n_1590);
 assign sub_1033_2_n_51 = ~(in1_119_10_ | ~n_1556);
 assign sub_1033_2_n_50 = ~(in1_119_13_ | ~n_1578);
 assign sub_1033_2_n_49 = ~(in1_119_18_ | ~n_1559);
 assign sub_1033_2_n_48 = ~(in1_119_7_ & ~n_1480);
 assign sub_1033_2_n_47 = ~(in1_119_7_ | ~n_1480);
 assign sub_1033_2_n_46 = ~(in1_119_11_ | ~n_1596);
 assign sub_1033_2_n_45 = ~(in1_119_17_ | ~n_1473);
 assign sub_1033_2_n_44 = ~(in1_119_1_ & ~n_1478);
 assign sub_1033_2_n_43 = ~(in1_119_21_ & ~n_1592);
 assign sub_1033_2_n_42 = ~(in1_119_15_ | ~n_1550);
 assign sub_1033_2_n_41 = ~(in1_119_12_ | ~n_1582);
 assign sub_1033_2_n_40 = ~(in1_119_21_ | ~n_1592);
 assign sub_1033_2_n_39 = ~(in1_119_13_ & ~n_1578);
 assign sub_1033_2_n_38 = ~(in1_119_4_ | ~n_1570);
 assign sub_1033_2_n_37 = ~(in1_119_16_ | ~n_1563);
 assign sub_1033_2_n_36 = ~(n_1544 & ~n_1402);
 assign sub_1033_2_n_35 = ~n_1544;
 assign sub_1033_2_n_34 = ~n_1587;
 assign in1_121_14_ = ~(sub_1033_2_n_152 ^ sub_1033_2_n_2);
 assign sub_1033_2_n_32 = (sub_1033_2_n_147 & sub_1033_2_n_126);
 assign sub_1033_2_n_31 = ~(sub_1033_2_n_112 | ~sub_1033_2_n_142);
 assign in1_121_23_ = (sub_1033_2_n_167 ^ sub_1033_2_n_99);
 assign sub_1033_2_n_29 = ~(sub_1033_2_n_93 | ~sub_1033_2_n_98);
 assign in1_121_22_ = (sub_1033_2_n_165 ^ sub_1033_2_n_3);
 assign in1_121_21_ = (sub_1033_2_n_164 ^ sub_1033_2_n_95);
 assign in1_121_11_ = (sub_1033_2_n_148 ^ sub_1033_2_n_94);
 assign in1_121_6_ = ~(sub_1033_2_n_138 ^ sub_1033_2_n_9);
 assign in1_121_19_ = (sub_1033_2_n_163 ^ sub_1033_2_n_91);
 assign in1_121_4_ = ~(sub_1033_2_n_130 ^ sub_1033_2_n_12);
 assign sub_1033_2_n_22 = ~(sub_1033_2_n_142 | ~sub_1033_2_n_87);
 assign in1_121_7_ = (sub_1033_2_n_143 ^ sub_1033_2_n_86);
 assign in1_121_3_ = (sub_1033_2_n_132 ^ sub_1033_2_n_13);
 assign in1_121_9_ = (sub_1033_2_n_145 ^ sub_1033_2_n_5);
 assign in1_121_15_ = (sub_1033_2_n_160 ^ sub_1033_2_n_85);
 assign in1_121_13_ = (sub_1033_2_n_151 ^ sub_1033_2_n_6);
 assign sub_1033_2_n_16 = ~(sub_1033_2_n_32 | ~sub_1033_2_n_84);
 assign in1_121_17_ = (sub_1033_2_n_156 ^ sub_1033_2_n_82);
 assign in1_121_10_ = ~(sub_1033_2_n_31 ^ sub_1033_2_n_8);
 assign sub_1033_2_n_13 = ~(sub_1033_2_n_72 | ~sub_1033_2_n_78);
 assign sub_1033_2_n_12 = ~(sub_1033_2_n_59 | ~sub_1033_2_n_73);
 assign sub_1033_2_n_11 = (sub_1033_2_n_72 | sub_1033_2_n_66);
 assign sub_1033_2_n_10 = ~(sub_1033_2_n_46 | ~sub_1033_2_n_70);
 assign sub_1033_2_n_9 = ~(sub_1033_2_n_68 | ~sub_1033_2_n_63);
 assign sub_1033_2_n_8 = ~(sub_1033_2_n_1 | ~sub_1033_2_n_61);
 assign sub_1033_2_n_7 = ~(sub_1033_2_n_38 | ~sub_1033_2_n_57);
 assign sub_1033_2_n_6 = ~(sub_1033_2_n_41 | ~sub_1033_2_n_54);
 assign sub_1033_2_n_5 = ~(sub_1033_2_n_0 | ~sub_1033_2_n_52);
 assign sub_1033_2_n_4 = ~(sub_1033_2_n_47 | ~sub_1033_2_n_48);
 assign sub_1033_2_n_3 = ~(sub_1033_2_n_40 | ~sub_1033_2_n_43);
 assign sub_1033_2_n_2 = ~(sub_1033_2_n_50 | ~sub_1033_2_n_39);
 assign sub_1033_2_n_1 = ~(in1_119_9_ | ~n_1552);
 assign sub_1033_2_n_0 = ~(in1_119_8_ | ~n_1590);
 assign sub_1054_2_n_167 = ~(sub_1054_2_n_42 & (sub_1054_2_n_166 | sub_1054_2_n_0));
 assign in1_124_24_ = (sub_1054_2_n_155 ^ in1_122_23_);
 assign sub_1054_2_n_164 = ~(sub_1054_2_n_61 & (sub_1054_2_n_157 | sub_1054_2_n_6));
 assign sub_1054_2_n_163 = ~(sub_1054_2_n_33 & (sub_1054_2_n_159 | sub_1054_2_n_4));
 assign sub_1054_2_n_162 = ~(sub_1054_2_n_34 & (sub_1054_2_n_158 | sub_1054_2_n_38));
 assign sub_1054_2_n_166 = ~(sub_1054_2_n_107 | (sub_1054_2_n_156 & sub_1054_2_n_75));
 assign in1_124_20_ = ~(sub_1054_2_n_156 ^ sub_1054_2_n_87);
 assign in1_124_13_ = (sub_1054_2_n_152 ^ sub_1054_2_n_71);
 assign sub_1054_2_n_157 = ~sub_1054_2_n_156;
 assign sub_1054_2_n_155 = ~(sub_1054_2_n_131 | ((sub_1054_2_n_144 & sub_1054_2_n_119) | (sub_1054_2_n_133
    & sub_1054_2_n_119)));
 assign sub_1054_2_n_154 = ~(sub_1054_2_n_32 & (sub_1054_2_n_149 | sub_1054_2_n_59));
 assign sub_1054_2_n_159 = ~(sub_1054_2_n_108 | (sub_1054_2_n_148 & sub_1054_2_n_102));
 assign sub_1054_2_n_158 = ~(sub_1054_2_n_109 | (sub_1054_2_n_147 & sub_1054_2_n_74));
 assign sub_1054_2_n_156 = ~(sub_1054_2_n_125 & (sub_1054_2_n_149 | sub_1054_2_n_115));
 assign in1_124_16_ = ~(sub_1054_2_n_149 ^ sub_1054_2_n_72);
 assign sub_1054_2_n_152 = ~(sub_1054_2_n_37 | (sub_1054_2_n_147 & sub_1054_2_n_51));
 assign sub_1054_2_n_151 = ~(sub_1054_2_n_53 & (sub_1054_2_n_23 | sub_1054_2_n_55));
 assign in1_124_7_ = (sub_1054_2_n_143 ^ sub_1054_2_n_88);
 assign sub_1054_2_n_148 = ~sub_1054_2_n_149;
 assign sub_1054_2_n_149 = ~(sub_1054_2_n_144 | sub_1054_2_n_133);
 assign sub_1054_2_n_147 = ~(sub_1054_2_n_124 & (sub_1054_2_n_141 | sub_1054_2_n_21));
 assign sub_1054_2_n_146 = ~(sub_1054_2_n_30 & (sub_1054_2_n_141 | sub_1054_2_n_35));
 assign in1_124_8_ = ~(sub_1054_2_n_141 ^ sub_1054_2_n_70);
 assign sub_1054_2_n_144 = ~(sub_1054_2_n_141 | sub_1054_2_n_120);
 assign sub_1054_2_n_143 = ~(sub_1054_2_n_58 & (sub_1054_2_n_140 | sub_1054_2_n_1));
 assign in1_124_5_ = ~(sub_1054_2_n_139 ^ sub_1054_2_n_90);
 assign sub_1054_2_n_141 = ~(sub_1054_2_n_123 | (sub_1054_2_n_137 & sub_1054_2_n_78));
 assign sub_1054_2_n_140 = ~(sub_1054_2_n_137 | sub_1054_2_n_110);
 assign sub_1054_2_n_139 = ~(sub_1054_2_n_41 & (sub_1054_2_n_134 | sub_1054_2_n_43));
 assign in1_124_3_ = (sub_1054_2_n_136 ^ sub_1054_2_n_91);
 assign sub_1054_2_n_137 = ~(sub_1054_2_n_134 | sub_1054_2_n_92);
 assign sub_1054_2_n_136 = ~(sub_1054_2_n_39 & (sub_1054_2_n_130 | sub_1054_2_n_54));
 assign in1_124_2_ = ~(sub_1054_2_n_130 ^ sub_1054_2_n_89);
 assign sub_1054_2_n_134 = ~(sub_1054_2_n_132 | sub_1054_2_n_112);
 assign sub_1054_2_n_133 = ~(sub_1054_2_n_127 & (sub_1054_2_n_124 | sub_1054_2_n_118));
 assign sub_1054_2_n_132 = ~(sub_1054_2_n_130 | sub_1054_2_n_8);
 assign sub_1054_2_n_131 = ~(sub_1054_2_n_24 & sub_1054_2_n_126);
 assign sub_1054_2_n_130 = ~(sub_1054_2_n_129 | sub_1054_2_n_113);
 assign sub_1054_2_n_129 = ~(sub_1054_2_n_122 & ~(sub_1054_2_n_49 & in1_122_0_));
 assign in1_124_1_ = (sub_1054_2_n_114 ^ sub_1054_2_n_49);
 assign sub_1054_2_n_127 = ~(sub_1054_2_n_103 | (sub_1054_2_n_109 & sub_1054_2_n_86));
 assign sub_1054_2_n_126 = ~(sub_1054_2_n_20 | sub_1054_2_n_105);
 assign sub_1054_2_n_125 = ~(sub_1054_2_n_106 | (sub_1054_2_n_108 & sub_1054_2_n_94));
 assign sub_1054_2_n_124 = ~(sub_1054_2_n_121 | sub_1054_2_n_111);
 assign sub_1054_2_n_123 = ~(sub_1054_2_n_104 & ~(sub_1054_2_n_110 & sub_1054_2_n_78));
 assign sub_1054_2_n_122 = ~(sub_1054_2_n_49 & ~n_1587);
 assign sub_1054_2_n_121 = ~(sub_1054_2_n_116 | sub_1054_2_n_100);
 assign sub_1054_2_n_120 = (sub_1054_2_n_21 | sub_1054_2_n_118);
 assign sub_1054_2_n_119 = ~(sub_1054_2_n_115 | sub_1054_2_n_117);
 assign sub_1054_2_n_113 = (sub_1054_2_n_28 & in1_122_0_);
 assign sub_1054_2_n_114 = (sub_1054_2_n_28 ^ in1_122_0_);
 assign sub_1054_2_n_112 = ~(sub_1054_2_n_65 & (sub_1054_2_n_39 | sub_1054_2_n_56));
 assign sub_1054_2_n_111 = ~(sub_1054_2_n_68 & (sub_1054_2_n_53 | sub_1054_2_n_7));
 assign sub_1054_2_n_118 = ~(sub_1054_2_n_74 & sub_1054_2_n_86);
 assign sub_1054_2_n_117 = ~(sub_1054_2_n_75 & sub_1054_2_n_99);
 assign sub_1054_2_n_116 = ~(sub_1054_2_n_64 | ~(sub_1054_2_n_30 | sub_1054_2_n_52));
 assign sub_1054_2_n_115 = ~(sub_1054_2_n_102 & sub_1054_2_n_94);
 assign sub_1054_2_n_106 = ~(sub_1054_2_n_46 & (sub_1054_2_n_33 | sub_1054_2_n_62));
 assign sub_1054_2_n_105 = ~(sub_1054_2_n_47 & (sub_1054_2_n_42 | sub_1054_2_n_2));
 assign sub_1054_2_n_104 = ~(sub_1054_2_n_66 | ~(sub_1054_2_n_58 | sub_1054_2_n_31));
 assign sub_1054_2_n_103 = ~(sub_1054_2_n_45 & (sub_1054_2_n_34 | sub_1054_2_n_63));
 assign sub_1054_2_n_110 = ~(sub_1054_2_n_44 & (sub_1054_2_n_41 | sub_1054_2_n_57));
 assign sub_1054_2_n_109 = ~(sub_1054_2_n_69 & (sub_1054_2_n_36 | sub_1054_2_n_60));
 assign sub_1054_2_n_108 = ~(sub_1054_2_n_48 & (sub_1054_2_n_32 | sub_1054_2_n_3));
 assign sub_1054_2_n_107 = ~(sub_1054_2_n_67 & (sub_1054_2_n_61 | sub_1054_2_n_5));
 assign sub_1054_2_n_92 = (sub_1054_2_n_43 | sub_1054_2_n_57);
 assign sub_1054_2_n_102 = ~(sub_1054_2_n_59 | sub_1054_2_n_3);
 assign sub_1054_2_n_101 = ~(sub_1054_2_n_1 | ~sub_1054_2_n_58);
 assign sub_1054_2_n_91 = ~(sub_1054_2_n_56 | ~sub_1054_2_n_65);
 assign sub_1054_2_n_90 = ~(sub_1054_2_n_44 & ~sub_1054_2_n_57);
 assign sub_1054_2_n_89 = ~(sub_1054_2_n_54 | ~sub_1054_2_n_39);
 assign sub_1054_2_n_100 = ~(sub_1054_2_n_40 & ~sub_1054_2_n_55);
 assign sub_1054_2_n_99 = ~(sub_1054_2_n_0 | sub_1054_2_n_2);
 assign sub_1054_2_n_98 = ~(sub_1054_2_n_2 | ~sub_1054_2_n_47);
 assign sub_1054_2_n_97 = ~(sub_1054_2_n_64 | sub_1054_2_n_52);
 assign sub_1054_2_n_96 = ~(sub_1054_2_n_0 | ~sub_1054_2_n_42);
 assign sub_1054_2_n_95 = ~(sub_1054_2_n_5 | ~sub_1054_2_n_67);
 assign sub_1054_2_n_88 = ~(sub_1054_2_n_66 | sub_1054_2_n_31);
 assign sub_1054_2_n_94 = ~(sub_1054_2_n_4 | sub_1054_2_n_62);
 assign sub_1054_2_n_87 = ~(sub_1054_2_n_61 & ~sub_1054_2_n_6);
 assign sub_1054_2_n_93 = ~(sub_1054_2_n_62 | ~sub_1054_2_n_46);
 assign in1_124_0_ = ~(sub_1054_2_n_49 & ~(sub_1054_2_n_29 & n_1598));
 assign sub_1054_2_n_86 = ~(sub_1054_2_n_38 | sub_1054_2_n_63);
 assign sub_1054_2_n_85 = ~(sub_1054_2_n_4 | ~sub_1054_2_n_33);
 assign sub_1054_2_n_84 = ~(sub_1054_2_n_43 | ~sub_1054_2_n_41);
 assign sub_1054_2_n_83 = ~(sub_1054_2_n_3 | ~sub_1054_2_n_48);
 assign sub_1054_2_n_72 = ~(sub_1054_2_n_59 | ~sub_1054_2_n_32);
 assign sub_1054_2_n_82 = ~(sub_1054_2_n_68 & sub_1054_2_n_40);
 assign sub_1054_2_n_81 = ~(sub_1054_2_n_38 | ~sub_1054_2_n_34);
 assign sub_1054_2_n_80 = ~(sub_1054_2_n_36 & sub_1054_2_n_51);
 assign sub_1054_2_n_79 = ~(sub_1054_2_n_35 | sub_1054_2_n_52);
 assign sub_1054_2_n_71 = ~(sub_1054_2_n_69 & ~sub_1054_2_n_60);
 assign sub_1054_2_n_78 = ~(sub_1054_2_n_1 | sub_1054_2_n_31);
 assign sub_1054_2_n_70 = ~(sub_1054_2_n_35 | ~sub_1054_2_n_30);
 assign sub_1054_2_n_77 = ~(sub_1054_2_n_63 | ~sub_1054_2_n_45);
 assign sub_1054_2_n_76 = ~(sub_1054_2_n_55 | ~sub_1054_2_n_53);
 assign sub_1054_2_n_75 = ~(sub_1054_2_n_6 | sub_1054_2_n_5);
 assign sub_1054_2_n_74 = ~(sub_1054_2_n_50 | sub_1054_2_n_60);
 assign sub_1054_2_n_51 = ~sub_1054_2_n_50;
 assign sub_1054_2_n_69 = ~(in1_122_12_ & ~n_1582);
 assign sub_1054_2_n_68 = ~(in1_122_10_ & ~n_1556);
 assign sub_1054_2_n_67 = ~(in1_122_20_ & ~n_1594);
 assign sub_1054_2_n_66 = ~(n_1528 | ~in1_122_6_);
 assign sub_1054_2_n_65 = ~(in1_122_2_ & ~n_1580);
 assign sub_1054_2_n_64 = ~(n_1590 | ~in1_122_8_);
 assign sub_1054_2_n_63 = ~(in1_122_14_ | ~n_1496);
 assign sub_1054_2_n_62 = ~(in1_122_18_ | ~n_1559);
 assign sub_1054_2_n_61 = ~(in1_122_19_ & ~n_1566);
 assign sub_1054_2_n_60 = ~(in1_122_12_ | ~n_1582);
 assign sub_1054_2_n_59 = ~(in1_122_15_ | ~n_1550);
 assign sub_1054_2_n_58 = ~(in1_122_5_ & ~n_1568);
 assign sub_1054_2_n_57 = ~(in1_122_4_ | ~n_1570);
 assign sub_1054_2_n_56 = ~(in1_122_2_ | ~n_1580);
 assign sub_1054_2_n_55 = ~(in1_122_9_ | ~n_1552);
 assign sub_1054_2_n_54 = ~(in1_122_1_ | ~n_1478);
 assign sub_1054_2_n_53 = ~(in1_122_9_ & ~n_1552);
 assign sub_1054_2_n_52 = ~(in1_122_8_ | ~n_1590);
 assign sub_1054_2_n_50 = ~(in1_122_11_ | ~n_1596);
 assign sub_1054_2_n_49 = ~(n_1544 & ~n_1598);
 assign sub_1054_2_n_40 = ~sub_1054_2_n_7;
 assign sub_1054_2_n_37 = ~sub_1054_2_n_36;
 assign sub_1054_2_n_48 = ~(in1_122_16_ & ~n_1563);
 assign sub_1054_2_n_47 = ~(in1_122_22_ & ~n_1404);
 assign sub_1054_2_n_46 = ~(in1_122_18_ & ~n_1559);
 assign sub_1054_2_n_45 = ~(in1_122_14_ & ~n_1496);
 assign sub_1054_2_n_44 = ~(in1_122_4_ & ~n_1570);
 assign sub_1054_2_n_43 = ~(in1_122_3_ | ~n_1536);
 assign sub_1054_2_n_42 = ~(in1_122_21_ & ~n_1592);
 assign sub_1054_2_n_41 = ~(in1_122_3_ & ~n_1536);
 assign sub_1054_2_n_39 = ~(in1_122_1_ & ~n_1478);
 assign sub_1054_2_n_38 = ~(in1_122_13_ | ~n_1578);
 assign sub_1054_2_n_36 = ~(in1_122_11_ & ~n_1596);
 assign sub_1054_2_n_35 = ~(in1_122_7_ | ~n_1480);
 assign sub_1054_2_n_34 = ~(in1_122_13_ & ~n_1578);
 assign sub_1054_2_n_33 = ~(in1_122_17_ & ~n_1473);
 assign sub_1054_2_n_32 = ~(in1_122_15_ & ~n_1550);
 assign sub_1054_2_n_31 = ~(in1_122_6_ | ~n_1528);
 assign sub_1054_2_n_30 = ~(in1_122_7_ & ~n_1480);
 assign sub_1054_2_n_29 = ~n_1544;
 assign sub_1054_2_n_28 = ~n_1587;
 assign in1_124_18_ = ~(sub_1054_2_n_159 ^ sub_1054_2_n_85);
 assign in1_124_14_ = ~(sub_1054_2_n_158 ^ sub_1054_2_n_81);
 assign in1_124_10_ = ~(sub_1054_2_n_23 ^ sub_1054_2_n_76);
 assign sub_1054_2_n_24 = (sub_1054_2_n_117 | sub_1054_2_n_125);
 assign sub_1054_2_n_23 = ~(sub_1054_2_n_10 | ~sub_1054_2_n_116);
 assign in1_124_6_ = ~(sub_1054_2_n_140 ^ sub_1054_2_n_101);
 assign sub_1054_2_n_21 = ~(sub_1054_2_n_79 & ~sub_1054_2_n_100);
 assign sub_1054_2_n_20 = (sub_1054_2_n_99 & sub_1054_2_n_107);
 assign in1_124_23_ = (sub_1054_2_n_167 ^ sub_1054_2_n_98);
 assign in1_124_9_ = (sub_1054_2_n_146 ^ sub_1054_2_n_97);
 assign in1_124_22_ = ~(sub_1054_2_n_166 ^ sub_1054_2_n_96);
 assign in1_124_21_ = (sub_1054_2_n_164 ^ sub_1054_2_n_95);
 assign in1_124_19_ = (sub_1054_2_n_163 ^ sub_1054_2_n_93);
 assign in1_124_4_ = ~(sub_1054_2_n_134 ^ sub_1054_2_n_84);
 assign in1_124_17_ = (sub_1054_2_n_154 ^ sub_1054_2_n_83);
 assign in1_124_11_ = ~(sub_1054_2_n_151 ^ sub_1054_2_n_82);
 assign in1_124_12_ = ~(sub_1054_2_n_147 ^ sub_1054_2_n_80);
 assign sub_1054_2_n_10 = ~(sub_1054_2_n_141 | ~sub_1054_2_n_79);
 assign in1_124_15_ = (sub_1054_2_n_162 ^ sub_1054_2_n_77);
 assign sub_1054_2_n_8 = (sub_1054_2_n_56 | sub_1054_2_n_54);
 assign sub_1054_2_n_7 = ~(in1_122_10_ | ~n_1556);
 assign sub_1054_2_n_6 = ~(in1_122_19_ | ~n_1566);
 assign sub_1054_2_n_5 = ~(in1_122_20_ | ~n_1594);
 assign sub_1054_2_n_4 = ~(in1_122_17_ | ~n_1473);
 assign sub_1054_2_n_3 = ~(in1_122_16_ | ~n_1563);
 assign sub_1054_2_n_2 = ~(in1_122_22_ | ~n_1404);
 assign sub_1054_2_n_1 = ~(in1_122_5_ | ~n_1568);
 assign sub_1054_2_n_0 = ~(in1_122_21_ | ~n_1592);
 assign in1_127_23_ = ~(sub_1075_2_n_183 ^ sub_1075_2_n_95);
 assign sub_1075_2_n_183 = ~(sub_1075_2_n_47 | (sub_1075_2_n_182 & sub_1075_2_n_43));
 assign sub_1075_2_n_182 = ~sub_1075_2_n_181;
 assign in1_127_24_ = ~(sub_1075_2_n_168 ^ in1_125_23_);
 assign sub_1075_2_n_179 = ~(sub_1075_2_n_172 | sub_1075_2_n_65);
 assign sub_1075_2_n_178 = ~(sub_1075_2_n_171 | sub_1075_2_n_33);
 assign sub_1075_2_n_177 = ~(sub_1075_2_n_35 | ~(sub_1075_2_n_22 | sub_1075_2_n_39));
 assign sub_1075_2_n_181 = ~(sub_1075_2_n_173 | sub_1075_2_n_113);
 assign in1_127_20_ = ~(sub_1075_2_n_169 ^ sub_1075_2_n_93);
 assign in1_127_14_ = ~(sub_1075_2_n_22 ^ sub_1075_2_n_78);
 assign in1_127_13_ = (sub_1075_2_n_165 ^ sub_1075_2_n_76);
 assign sub_1075_2_n_173 = ~(sub_1075_2_n_169 | sub_1075_2_n_82);
 assign sub_1075_2_n_172 = ~(sub_1075_2_n_169 | sub_1075_2_n_60);
 assign sub_1075_2_n_171 = ~(sub_1075_2_n_170 | sub_1075_2_n_32);
 assign sub_1075_2_n_168 = ~(sub_1075_2_n_160 & sub_1075_2_n_144);
 assign sub_1075_2_n_167 = ~(sub_1075_2_n_163 | sub_1075_2_n_31);
 assign sub_1075_2_n_170 = ~(sub_1075_2_n_17 | sub_1075_2_n_114);
 assign sub_1075_2_n_169 = ~(sub_1075_2_n_131 | ~(sub_1075_2_n_159 | sub_1075_2_n_121));
 assign in1_127_12_ = ~(sub_1075_2_n_158 ^ sub_1075_2_n_77);
 assign sub_1075_2_n_165 = ~(sub_1075_2_n_38 | ~(sub_1075_2_n_158 | sub_1075_2_n_54));
 assign sub_1075_2_n_164 = ~(sub_1075_2_n_161 | sub_1075_2_n_56);
 assign sub_1075_2_n_163 = ~(sub_1075_2_n_159 | sub_1075_2_n_2);
 assign sub_1075_2_n_162 = ~(sub_1075_2_n_158 | sub_1075_2_n_8);
 assign sub_1075_2_n_161 = ~(sub_1075_2_n_157 | sub_1075_2_n_58);
 assign sub_1075_2_n_160 = ~(sub_1075_2_n_137 | (sub_1075_2_n_153 & sub_1075_2_n_23));
 assign sub_1075_2_n_159 = ~(sub_1075_2_n_153 | sub_1075_2_n_139);
 assign sub_1075_2_n_158 = ~(sub_1075_2_n_130 | ~(sub_1075_2_n_149 | sub_1075_2_n_123));
 assign sub_1075_2_n_157 = ~(sub_1075_2_n_154 | sub_1075_2_n_124);
 assign sub_1075_2_n_156 = ~(sub_1075_2_n_28 | ~(sub_1075_2_n_149 | sub_1075_2_n_36));
 assign in1_127_8_ = ~(sub_1075_2_n_149 ^ sub_1075_2_n_75);
 assign sub_1075_2_n_154 = ~(sub_1075_2_n_149 | sub_1075_2_n_87);
 assign sub_1075_2_n_153 = ~(sub_1075_2_n_149 | sub_1075_2_n_126);
 assign sub_1075_2_n_152 = ~(sub_1075_2_n_62 | (sub_1075_2_n_24 & sub_1075_2_n_1));
 assign in1_127_6_ = ~(sub_1075_2_n_24 ^ sub_1075_2_n_94);
 assign in1_127_5_ = ~(sub_1075_2_n_148 ^ sub_1075_2_n_97);
 assign sub_1075_2_n_149 = ~(sub_1075_2_n_129 | (sub_1075_2_n_145 & sub_1075_2_n_86));
 assign sub_1075_2_n_148 = ~(sub_1075_2_n_45 | (sub_1075_2_n_141 & sub_1075_2_n_5));
 assign in1_127_4_ = ~(sub_1075_2_n_141 ^ sub_1075_2_n_79);
 assign in1_127_3_ = ~(sub_1075_2_n_143 ^ sub_1075_2_n_98);
 assign sub_1075_2_n_145 = ~(sub_1075_2_n_140 | sub_1075_2_n_7);
 assign sub_1075_2_n_144 = ~(sub_1075_2_n_139 & sub_1075_2_n_23);
 assign sub_1075_2_n_143 = ~(sub_1075_2_n_40 & (sub_1075_2_n_136 | sub_1075_2_n_57));
 assign in1_127_2_ = ~(sub_1075_2_n_136 ^ sub_1075_2_n_96);
 assign sub_1075_2_n_141 = ~sub_1075_2_n_140;
 assign sub_1075_2_n_140 = ~(sub_1075_2_n_138 | sub_1075_2_n_118);
 assign sub_1075_2_n_139 = ~(sub_1075_2_n_133 & ~(sub_1075_2_n_130 & sub_1075_2_n_125));
 assign sub_1075_2_n_138 = ~(sub_1075_2_n_136 | sub_1075_2_n_6);
 assign sub_1075_2_n_137 = ~(sub_1075_2_n_132 & ~(sub_1075_2_n_131 & sub_1075_2_n_20));
 assign sub_1075_2_n_136 = ~(sub_1075_2_n_135 | sub_1075_2_n_119);
 assign sub_1075_2_n_135 = ~(sub_1075_2_n_128 & ~(sub_1075_2_n_53 & in1_125_0_));
 assign in1_127_1_ = (sub_1075_2_n_120 ^ sub_1075_2_n_53);
 assign sub_1075_2_n_133 = ~(sub_1075_2_n_127 | sub_1075_2_n_109);
 assign sub_1075_2_n_132 = ~(sub_1075_2_n_111 | (sub_1075_2_n_113 & sub_1075_2_n_106));
 assign sub_1075_2_n_131 = ~(sub_1075_2_n_112 & ~(sub_1075_2_n_114 & sub_1075_2_n_102));
 assign sub_1075_2_n_130 = ~(sub_1075_2_n_117 & ~(sub_1075_2_n_124 & sub_1075_2_n_107));
 assign sub_1075_2_n_129 = ~(sub_1075_2_n_110 & (sub_1075_2_n_116 | sub_1075_2_n_85));
 assign sub_1075_2_n_128 = ~(sub_1075_2_n_53 & ~n_1587);
 assign sub_1075_2_n_127 = ~(sub_1075_2_n_115 | sub_1075_2_n_92);
 assign sub_1075_2_n_126 = ~(sub_1075_2_n_122 & sub_1075_2_n_125);
 assign sub_1075_2_n_123 = ~sub_1075_2_n_122;
 assign sub_1075_2_n_119 = (sub_1075_2_n_25 & in1_125_0_);
 assign sub_1075_2_n_120 = (sub_1075_2_n_25 ^ in1_125_0_);
 assign sub_1075_2_n_118 = ~(sub_1075_2_n_70 & (sub_1075_2_n_40 | sub_1075_2_n_59));
 assign sub_1075_2_n_117 = ~(sub_1075_2_n_73 | (sub_1075_2_n_56 & sub_1075_2_n_42));
 assign sub_1075_2_n_125 = ~(sub_1075_2_n_8 | sub_1075_2_n_92);
 assign sub_1075_2_n_124 = ~(sub_1075_2_n_69 & (sub_1075_2_n_27 | sub_1075_2_n_55));
 assign sub_1075_2_n_122 = ~(sub_1075_2_n_87 | ~sub_1075_2_n_107);
 assign sub_1075_2_n_121 = ~(sub_1075_2_n_103 & sub_1075_2_n_102);
 assign sub_1075_2_n_112 = ~(sub_1075_2_n_50 | (sub_1075_2_n_33 & sub_1075_2_n_67));
 assign sub_1075_2_n_111 = ~(sub_1075_2_n_51 & (sub_1075_2_n_46 | sub_1075_2_n_3));
 assign sub_1075_2_n_110 = ~(sub_1075_2_n_81 | sub_1075_2_n_71);
 assign sub_1075_2_n_109 = ~(sub_1075_2_n_49 & ~(sub_1075_2_n_35 & sub_1075_2_n_68));
 assign sub_1075_2_n_116 = ~(sub_1075_2_n_99 | sub_1075_2_n_48);
 assign sub_1075_2_n_115 = ~(sub_1075_2_n_74 | ~(sub_1075_2_n_37 | sub_1075_2_n_63));
 assign sub_1075_2_n_114 = ~(sub_1075_2_n_52 & (sub_1075_2_n_30 | sub_1075_2_n_4));
 assign sub_1075_2_n_113 = ~(sub_1075_2_n_72 & (sub_1075_2_n_64 | sub_1075_2_n_34));
 assign sub_1075_2_n_99 = ~(sub_1075_2_n_44 | sub_1075_2_n_61);
 assign sub_1075_2_n_108 = ~(sub_1075_2_n_55 | ~sub_1075_2_n_69);
 assign sub_1075_2_n_98 = ~(sub_1075_2_n_70 & ~sub_1075_2_n_59);
 assign sub_1075_2_n_97 = ~(sub_1075_2_n_48 | sub_1075_2_n_61);
 assign sub_1075_2_n_96 = ~(sub_1075_2_n_57 | ~sub_1075_2_n_40);
 assign sub_1075_2_n_107 = ~(sub_1075_2_n_58 | sub_1075_2_n_41);
 assign sub_1075_2_n_106 = ~(sub_1075_2_n_0 | sub_1075_2_n_3);
 assign sub_1075_2_n_95 = ~(sub_1075_2_n_3 | ~sub_1075_2_n_51);
 assign sub_1075_2_n_94 = ~(sub_1075_2_n_1 & ~sub_1075_2_n_62);
 assign sub_1075_2_n_105 = ~(sub_1075_2_n_46 & sub_1075_2_n_43);
 assign sub_1075_2_n_104 = ~(sub_1075_2_n_34 | ~sub_1075_2_n_72);
 assign sub_1075_2_n_103 = ~(sub_1075_2_n_2 | sub_1075_2_n_4);
 assign sub_1075_2_n_102 = ~(sub_1075_2_n_32 | sub_1075_2_n_66);
 assign sub_1075_2_n_93 = ~(sub_1075_2_n_65 | sub_1075_2_n_60);
 assign sub_1075_2_n_101 = ~(sub_1075_2_n_50 | ~sub_1075_2_n_67);
 assign sub_1075_2_n_100 = ~(sub_1075_2_n_71 | sub_1075_2_n_29);
 assign sub_1075_2_n_86 = ~sub_1075_2_n_85;
 assign sub_1075_2_n_81 = ~(sub_1075_2_n_29 | ~sub_1075_2_n_62);
 assign in1_127_0_ = ~(sub_1075_2_n_53 & ~(sub_1075_2_n_26 & n_1576));
 assign sub_1075_2_n_92 = ~(sub_1075_2_n_68 & ~sub_1075_2_n_39);
 assign sub_1075_2_n_91 = ~(sub_1075_2_n_33 | sub_1075_2_n_32);
 assign sub_1075_2_n_79 = ~(sub_1075_2_n_44 & sub_1075_2_n_5);
 assign sub_1075_2_n_90 = ~(sub_1075_2_n_4 | ~sub_1075_2_n_52);
 assign sub_1075_2_n_89 = ~(sub_1075_2_n_31 | sub_1075_2_n_2);
 assign sub_1075_2_n_88 = ~(sub_1075_2_n_73 | sub_1075_2_n_41);
 assign sub_1075_2_n_78 = ~(sub_1075_2_n_35 | sub_1075_2_n_39);
 assign sub_1075_2_n_77 = ~(sub_1075_2_n_38 | sub_1075_2_n_54);
 assign sub_1075_2_n_87 = (sub_1075_2_n_36 | sub_1075_2_n_55);
 assign sub_1075_2_n_76 = (sub_1075_2_n_74 | sub_1075_2_n_63);
 assign sub_1075_2_n_85 = ~(sub_1075_2_n_1 & ~sub_1075_2_n_29);
 assign sub_1075_2_n_75 = ~(sub_1075_2_n_28 | sub_1075_2_n_36);
 assign sub_1075_2_n_84 = ~(sub_1075_2_n_49 & sub_1075_2_n_68);
 assign sub_1075_2_n_83 = ~(sub_1075_2_n_56 | sub_1075_2_n_58);
 assign sub_1075_2_n_82 = (sub_1075_2_n_60 | sub_1075_2_n_34);
 assign sub_1075_2_n_67 = ~sub_1075_2_n_66;
 assign sub_1075_2_n_65 = ~sub_1075_2_n_64;
 assign sub_1075_2_n_74 = ~(n_1582 | ~in1_125_12_);
 assign sub_1075_2_n_73 = ~(n_1556 | ~in1_125_10_);
 assign sub_1075_2_n_72 = ~(in1_125_20_ & ~n_1594);
 assign sub_1075_2_n_71 = ~(n_1528 | ~in1_125_6_);
 assign sub_1075_2_n_70 = ~(in1_125_2_ & ~n_1580);
 assign sub_1075_2_n_69 = ~(in1_125_8_ & ~n_1590);
 assign sub_1075_2_n_68 = ~(n_1496 & ~in1_125_14_);
 assign sub_1075_2_n_66 = ~(in1_125_18_ | ~n_1559);
 assign sub_1075_2_n_64 = ~(in1_125_19_ & ~n_1566);
 assign sub_1075_2_n_63 = ~(in1_125_12_ | ~n_1582);
 assign sub_1075_2_n_62 = ~(n_1568 | ~in1_125_5_);
 assign sub_1075_2_n_61 = ~(in1_125_4_ | ~n_1570);
 assign sub_1075_2_n_60 = ~(in1_125_19_ | ~n_1566);
 assign sub_1075_2_n_59 = ~(in1_125_2_ | ~n_1580);
 assign sub_1075_2_n_58 = ~(in1_125_9_ | ~n_1552);
 assign sub_1075_2_n_57 = ~(in1_125_1_ | ~n_1478);
 assign sub_1075_2_n_56 = ~(n_1552 | ~in1_125_9_);
 assign sub_1075_2_n_55 = ~(in1_125_8_ | ~n_1590);
 assign sub_1075_2_n_54 = ~(in1_125_11_ | ~n_1596);
 assign sub_1075_2_n_53 = ~(n_1544 & ~n_1576);
 assign sub_1075_2_n_47 = ~sub_1075_2_n_46;
 assign sub_1075_2_n_45 = ~sub_1075_2_n_44;
 assign sub_1075_2_n_43 = ~sub_1075_2_n_0;
 assign sub_1075_2_n_42 = ~sub_1075_2_n_41;
 assign sub_1075_2_n_38 = ~sub_1075_2_n_37;
 assign sub_1075_2_n_31 = ~sub_1075_2_n_30;
 assign sub_1075_2_n_28 = ~sub_1075_2_n_27;
 assign sub_1075_2_n_52 = ~(in1_125_16_ & ~n_1563);
 assign sub_1075_2_n_51 = ~(in1_125_22_ & ~n_1404);
 assign sub_1075_2_n_50 = ~(n_1559 | ~in1_125_18_);
 assign sub_1075_2_n_49 = ~(in1_125_14_ & ~n_1496);
 assign sub_1075_2_n_48 = ~(n_1570 | ~in1_125_4_);
 assign sub_1075_2_n_46 = ~(in1_125_21_ & ~n_1592);
 assign sub_1075_2_n_44 = ~(in1_125_3_ & ~n_1536);
 assign sub_1075_2_n_41 = ~(in1_125_10_ | ~n_1556);
 assign sub_1075_2_n_40 = ~(in1_125_1_ & ~n_1478);
 assign sub_1075_2_n_39 = ~(in1_125_13_ | ~n_1578);
 assign sub_1075_2_n_37 = ~(in1_125_11_ & ~n_1596);
 assign sub_1075_2_n_36 = ~(in1_125_7_ | ~n_1480);
 assign sub_1075_2_n_35 = ~(n_1578 | ~in1_125_13_);
 assign sub_1075_2_n_34 = ~(in1_125_20_ | ~n_1594);
 assign sub_1075_2_n_33 = ~(n_1473 | ~in1_125_17_);
 assign sub_1075_2_n_32 = ~(in1_125_17_ | ~n_1473);
 assign sub_1075_2_n_30 = ~(in1_125_15_ & ~n_1550);
 assign sub_1075_2_n_29 = ~(in1_125_6_ | ~n_1528);
 assign sub_1075_2_n_27 = ~(in1_125_7_ & ~n_1480);
 assign sub_1075_2_n_26 = ~n_1544;
 assign sub_1075_2_n_25 = ~n_1587;
 assign sub_1075_2_n_24 = ~(sub_1075_2_n_116 & ~sub_1075_2_n_145);
 assign sub_1075_2_n_23 = ~(sub_1075_2_n_121 | ~sub_1075_2_n_20);
 assign sub_1075_2_n_22 = ~(sub_1075_2_n_162 | ~sub_1075_2_n_115);
 assign in1_127_9_ = ~(sub_1075_2_n_156 ^ sub_1075_2_n_108);
 assign sub_1075_2_n_20 = ~(sub_1075_2_n_82 | ~sub_1075_2_n_106);
 assign in1_127_22_ = (sub_1075_2_n_181 ^ sub_1075_2_n_105);
 assign in1_127_21_ = ~(sub_1075_2_n_179 ^ sub_1075_2_n_104);
 assign sub_1075_2_n_17 = ~(sub_1075_2_n_159 | ~sub_1075_2_n_103);
 assign in1_127_19_ = ~(sub_1075_2_n_178 ^ sub_1075_2_n_101);
 assign in1_127_7_ = ~(sub_1075_2_n_152 ^ sub_1075_2_n_100);
 assign in1_127_18_ = ~(sub_1075_2_n_170 ^ sub_1075_2_n_91);
 assign in1_127_17_ = ~(sub_1075_2_n_167 ^ sub_1075_2_n_90);
 assign in1_127_16_ = ~(sub_1075_2_n_159 ^ sub_1075_2_n_89);
 assign in1_127_11_ = ~(sub_1075_2_n_164 ^ sub_1075_2_n_88);
 assign in1_127_15_ = (sub_1075_2_n_177 ^ sub_1075_2_n_84);
 assign in1_127_10_ = ~(sub_1075_2_n_157 ^ sub_1075_2_n_83);
 assign sub_1075_2_n_8 = (sub_1075_2_n_63 | sub_1075_2_n_54);
 assign sub_1075_2_n_7 = ~(sub_1075_2_n_5 & ~sub_1075_2_n_61);
 assign sub_1075_2_n_6 = (sub_1075_2_n_59 | sub_1075_2_n_57);
 assign sub_1075_2_n_5 = ~(n_1536 & ~in1_125_3_);
 assign sub_1075_2_n_4 = ~(in1_125_16_ | ~n_1563);
 assign sub_1075_2_n_3 = ~(in1_125_22_ | ~n_1404);
 assign sub_1075_2_n_2 = ~(in1_125_15_ | ~n_1550);
 assign sub_1075_2_n_1 = ~(n_1568 & ~in1_125_5_);
 assign sub_1075_2_n_0 = ~(in1_125_21_ | ~n_1592);
 assign in1_130_23_ = ~(sub_1096_2_n_169 ^ sub_1096_2_n_79);
 assign sub_1096_2_n_169 = ~(sub_1096_2_n_16 & (sub_1096_2_n_166 | sub_1096_2_n_37));
 assign in1_130_21_ = ~(sub_1096_2_n_165 ^ sub_1096_2_n_76);
 assign in1_130_19_ = ~(sub_1096_2_n_164 ^ sub_1096_2_n_73);
 assign sub_1096_2_n_166 = ~(sub_1096_2_n_95 | (sub_1096_2_n_153 & sub_1096_2_n_83));
 assign sub_1096_2_n_165 = ~(sub_1096_2_n_15 & (sub_1096_2_n_152 | sub_1096_2_n_46));
 assign sub_1096_2_n_164 = ~(sub_1096_2_n_27 & (sub_1096_2_n_154 | sub_1096_2_n_41));
 assign sub_1096_2_n_163 = ~(sub_1096_2_n_48 & (sub_1096_2_n_155 | sub_1096_2_n_2));
 assign in1_130_20_ = ~(sub_1096_2_n_153 ^ sub_1096_2_n_75);
 assign in1_130_18_ = ~(sub_1096_2_n_154 ^ sub_1096_2_n_62);
 assign in1_130_17_ = ~(sub_1096_2_n_149 ^ sub_1096_2_n_65);
 assign in1_130_14_ = ~(sub_1096_2_n_155 ^ sub_1096_2_n_60);
 assign in1_130_13_ = ~(sub_1096_2_n_144 ^ sub_1096_2_n_59);
 assign in1_130_11_ = ~(sub_1096_2_n_143 ^ sub_1096_2_n_64);
 assign in1_130_24_ = (sub_1096_2_n_151 | sub_1096_2_n_150);
 assign sub_1096_2_n_153 = ~sub_1096_2_n_152;
 assign sub_1096_2_n_151 = ~(sub_1096_2_n_141 | in1_128_23_);
 assign sub_1096_2_n_150 = ~(sub_1096_2_n_140 | ~in1_128_23_);
 assign sub_1096_2_n_149 = ~(sub_1096_2_n_28 & (sub_1096_2_n_8 | sub_1096_2_n_19));
 assign sub_1096_2_n_155 = ~(sub_1096_2_n_96 | (sub_1096_2_n_137 & sub_1096_2_n_84));
 assign sub_1096_2_n_154 = ~(sub_1096_2_n_4 | sub_1096_2_n_94);
 assign sub_1096_2_n_152 = ~(sub_1096_2_n_142 | sub_1096_2_n_108);
 assign in1_130_10_ = ~(sub_1096_2_n_135 ^ sub_1096_2_n_57);
 assign in1_130_12_ = ~(sub_1096_2_n_137 ^ sub_1096_2_n_56);
 assign in1_130_16_ = ~(sub_1096_2_n_8 ^ sub_1096_2_n_81);
 assign in1_130_9_ = ~(sub_1096_2_n_134 ^ sub_1096_2_n_78);
 assign sub_1096_2_n_144 = ~(sub_1096_2_n_45 & ~(sub_1096_2_n_137 & sub_1096_2_n_39));
 assign sub_1096_2_n_143 = ~(sub_1096_2_n_40 & (sub_1096_2_n_136 | sub_1096_2_n_20));
 assign sub_1096_2_n_142 = ~(sub_1096_2_n_8 | sub_1096_2_n_101);
 assign sub_1096_2_n_141 = ~sub_1096_2_n_140;
 assign sub_1096_2_n_140 = ~(sub_1096_2_n_138 | ~sub_1096_2_n_120);
 assign in1_130_7_ = ~(sub_1096_2_n_132 ^ sub_1096_2_n_61);
 assign sub_1096_2_n_138 = ~(sub_1096_2_n_131 | sub_1096_2_n_105);
 assign sub_1096_2_n_137 = ~(sub_1096_2_n_111 & (sub_1096_2_n_128 | sub_1096_2_n_6));
 assign sub_1096_2_n_136 = ~sub_1096_2_n_135;
 assign sub_1096_2_n_135 = ~(sub_1096_2_n_93 & (sub_1096_2_n_128 | sub_1096_2_n_71));
 assign sub_1096_2_n_134 = ~(sub_1096_2_n_21 & (sub_1096_2_n_128 | sub_1096_2_n_43));
 assign in1_130_8_ = ~(sub_1096_2_n_128 ^ sub_1096_2_n_80);
 assign sub_1096_2_n_132 = ~(sub_1096_2_n_42 & (sub_1096_2_n_125 | sub_1096_2_n_0));
 assign sub_1096_2_n_131 = ~(sub_1096_2_n_127 & sub_1096_2_n_106);
 assign in1_130_6_ = ~(sub_1096_2_n_125 ^ sub_1096_2_n_77);
 assign in1_130_5_ = ~(sub_1096_2_n_124 ^ sub_1096_2_n_58);
 assign sub_1096_2_n_128 = ~sub_1096_2_n_127;
 assign sub_1096_2_n_127 = ~(sub_1096_2_n_126 & sub_1096_2_n_110);
 assign sub_1096_2_n_126 = ~(sub_1096_2_n_121 & sub_1096_2_n_89);
 assign sub_1096_2_n_125 = ~(sub_1096_2_n_121 | sub_1096_2_n_97);
 assign sub_1096_2_n_124 = ~(sub_1096_2_n_22 & (sub_1096_2_n_116 | sub_1096_2_n_25));
 assign in1_130_4_ = ~(sub_1096_2_n_116 ^ sub_1096_2_n_55);
 assign in1_130_3_ = ~(sub_1096_2_n_118 ^ sub_1096_2_n_63);
 assign sub_1096_2_n_121 = ~(sub_1096_2_n_116 | sub_1096_2_n_82);
 assign sub_1096_2_n_120 = ~(sub_1096_2_n_119 | sub_1096_2_n_114);
 assign sub_1096_2_n_119 = ~(sub_1096_2_n_115 | sub_1096_2_n_105);
 assign sub_1096_2_n_118 = ~(sub_1096_2_n_13 | (sub_1096_2_n_113 & sub_1096_2_n_18));
 assign in1_130_2_ = ~(sub_1096_2_n_113 ^ sub_1096_2_n_74);
 assign sub_1096_2_n_116 = ~(sub_1096_2_n_91 | (sub_1096_2_n_113 & sub_1096_2_n_67));
 assign sub_1096_2_n_115 = ~(sub_1096_2_n_109 | ~(sub_1096_2_n_111 | sub_1096_2_n_103));
 assign sub_1096_2_n_114 = ~(sub_1096_2_n_107 & ~(sub_1096_2_n_108 & sub_1096_2_n_102));
 assign sub_1096_2_n_113 = ((sub_1096_2_n_11 & in1_128_0_) | ((in1_128_0_ & sub_1096_2_n_10) | (sub_1096_2_n_10
    & sub_1096_2_n_11)));
 assign in1_130_1_ = (in1_128_0_ ^ (sub_1096_2_n_10 ^ sub_1096_2_n_11));
 assign sub_1096_2_n_111 = ~(sub_1096_2_n_92 | ~(sub_1096_2_n_93 | sub_1096_2_n_72));
 assign sub_1096_2_n_110 = ~(sub_1096_2_n_99 | (sub_1096_2_n_97 & sub_1096_2_n_89));
 assign sub_1096_2_n_109 = ~(sub_1096_2_n_100 & ~(sub_1096_2_n_96 & sub_1096_2_n_88));
 assign sub_1096_2_n_108 = ~(sub_1096_2_n_98 & ~(sub_1096_2_n_94 & sub_1096_2_n_85));
 assign sub_1096_2_n_107 = ~(sub_1096_2_n_104 | sub_1096_2_n_90);
 assign sub_1096_2_n_106 = ~(sub_1096_2_n_6 | sub_1096_2_n_103);
 assign sub_1096_2_n_105 = ~(sub_1096_2_n_102 & ~sub_1096_2_n_101);
 assign sub_1096_2_n_104 = ~(sub_1096_2_n_87 | ~sub_1096_2_n_95);
 assign sub_1096_2_n_100 = ~(sub_1096_2_n_32 | ~(sub_1096_2_n_48 | sub_1096_2_n_24));
 assign sub_1096_2_n_99 = ~(sub_1096_2_n_34 & (sub_1096_2_n_42 | sub_1096_2_n_44));
 assign sub_1096_2_n_98 = ~(sub_1096_2_n_53 | ~(sub_1096_2_n_27 | sub_1096_2_n_14));
 assign sub_1096_2_n_103 = ~(sub_1096_2_n_84 & sub_1096_2_n_88);
 assign sub_1096_2_n_102 = ~(sub_1096_2_n_87 | ~sub_1096_2_n_83);
 assign sub_1096_2_n_101 = ~(sub_1096_2_n_68 & sub_1096_2_n_85);
 assign sub_1096_2_n_92 = ~(sub_1096_2_n_52 & (sub_1096_2_n_40 | sub_1096_2_n_26));
 assign sub_1096_2_n_91 = ~(sub_1096_2_n_54 & (sub_1096_2_n_12 | sub_1096_2_n_3));
 assign sub_1096_2_n_90 = ~(sub_1096_2_n_31 & (sub_1096_2_n_16 | sub_1096_2_n_47));
 assign sub_1096_2_n_97 = ~(sub_1096_2_n_30 & (sub_1096_2_n_22 | sub_1096_2_n_23));
 assign sub_1096_2_n_96 = ~(sub_1096_2_n_51 & (sub_1096_2_n_45 | sub_1096_2_n_29));
 assign sub_1096_2_n_95 = ~(sub_1096_2_n_33 & (sub_1096_2_n_15 | sub_1096_2_n_35));
 assign sub_1096_2_n_94 = ~(sub_1096_2_n_49 & (sub_1096_2_n_28 | sub_1096_2_n_1));
 assign sub_1096_2_n_93 = ~(sub_1096_2_n_50 | ~(sub_1096_2_n_21 | sub_1096_2_n_36));
 assign sub_1096_2_n_82 = (sub_1096_2_n_25 | sub_1096_2_n_23);
 assign sub_1096_2_n_81 = ~(sub_1096_2_n_19 | ~sub_1096_2_n_28);
 assign sub_1096_2_n_80 = ~(sub_1096_2_n_43 | ~sub_1096_2_n_21);
 assign sub_1096_2_n_79 = ~(sub_1096_2_n_31 & ~sub_1096_2_n_47);
 assign sub_1096_2_n_89 = ~(sub_1096_2_n_0 | sub_1096_2_n_44);
 assign sub_1096_2_n_78 = (sub_1096_2_n_50 | sub_1096_2_n_36);
 assign sub_1096_2_n_88 = ~(sub_1096_2_n_2 | sub_1096_2_n_24);
 assign sub_1096_2_n_77 = ~(sub_1096_2_n_0 | ~sub_1096_2_n_42);
 assign sub_1096_2_n_87 = (sub_1096_2_n_37 | sub_1096_2_n_47);
 assign sub_1096_2_n_86 = ~(sub_1096_2_n_37 | ~sub_1096_2_n_16);
 assign sub_1096_2_n_76 = ~(sub_1096_2_n_33 & ~sub_1096_2_n_35);
 assign sub_1096_2_n_85 = ~(sub_1096_2_n_41 | sub_1096_2_n_14);
 assign sub_1096_2_n_84 = ~(sub_1096_2_n_38 | sub_1096_2_n_29);
 assign sub_1096_2_n_75 = ~(sub_1096_2_n_15 & ~sub_1096_2_n_46);
 assign sub_1096_2_n_74 = ~(sub_1096_2_n_12 & sub_1096_2_n_18);
 assign sub_1096_2_n_73 = (sub_1096_2_n_53 | sub_1096_2_n_14);
 assign sub_1096_2_n_83 = ~(sub_1096_2_n_46 | sub_1096_2_n_35);
 assign sub_1096_2_n_71 = ~sub_1096_2_n_70;
 assign sub_1096_2_n_67 = ~(sub_1096_2_n_17 | sub_1096_2_n_3);
 assign in1_130_0_ = ~(sub_1096_2_n_11 & ~(sub_1096_2_n_9 & n_1574));
 assign sub_1096_2_n_65 = ~(sub_1096_2_n_49 & ~sub_1096_2_n_1);
 assign sub_1096_2_n_64 = ~(sub_1096_2_n_52 & ~sub_1096_2_n_26);
 assign sub_1096_2_n_72 = (sub_1096_2_n_20 | sub_1096_2_n_26);
 assign sub_1096_2_n_70 = ~(sub_1096_2_n_43 | sub_1096_2_n_36);
 assign sub_1096_2_n_63 = ~(sub_1096_2_n_3 | ~sub_1096_2_n_54);
 assign sub_1096_2_n_62 = ~(sub_1096_2_n_41 | ~sub_1096_2_n_27);
 assign sub_1096_2_n_69 = ~(sub_1096_2_n_32 | sub_1096_2_n_24);
 assign sub_1096_2_n_61 = ~(sub_1096_2_n_34 & ~sub_1096_2_n_44);
 assign sub_1096_2_n_60 = ~(sub_1096_2_n_2 | ~sub_1096_2_n_48);
 assign sub_1096_2_n_59 = ~(sub_1096_2_n_51 & ~sub_1096_2_n_29);
 assign sub_1096_2_n_58 = ~(sub_1096_2_n_30 & ~sub_1096_2_n_23);
 assign sub_1096_2_n_68 = ~(sub_1096_2_n_19 | sub_1096_2_n_1);
 assign sub_1096_2_n_57 = ~(sub_1096_2_n_40 & ~sub_1096_2_n_20);
 assign sub_1096_2_n_56 = ~(sub_1096_2_n_45 & sub_1096_2_n_39);
 assign sub_1096_2_n_55 = ~(sub_1096_2_n_25 | ~sub_1096_2_n_22);
 assign sub_1096_2_n_39 = ~sub_1096_2_n_38;
 assign sub_1096_2_n_54 = ~(in1_128_2_ & ~n_1580);
 assign sub_1096_2_n_53 = ~(n_1559 | ~in1_128_18_);
 assign sub_1096_2_n_52 = ~(in1_128_10_ & ~n_1556);
 assign sub_1096_2_n_51 = ~(in1_128_12_ & ~n_1582);
 assign sub_1096_2_n_50 = ~(n_1590 | ~in1_128_8_);
 assign sub_1096_2_n_49 = ~(in1_128_16_ & ~n_1563);
 assign sub_1096_2_n_48 = ~(in1_128_13_ & ~n_1578);
 assign sub_1096_2_n_47 = ~(in1_128_22_ | ~n_1404);
 assign sub_1096_2_n_46 = ~(in1_128_19_ | ~n_1566);
 assign sub_1096_2_n_45 = ~(in1_128_11_ & ~n_1596);
 assign sub_1096_2_n_44 = ~(in1_128_6_ | ~n_1528);
 assign sub_1096_2_n_43 = ~(in1_128_7_ | ~n_1480);
 assign sub_1096_2_n_42 = ~(in1_128_5_ & ~n_1568);
 assign sub_1096_2_n_41 = ~(in1_128_17_ | ~n_1473);
 assign sub_1096_2_n_40 = ~(in1_128_9_ & ~n_1552);
 assign sub_1096_2_n_38 = ~(in1_128_11_ | ~n_1596);
 assign sub_1096_2_n_37 = ~(in1_128_21_ | ~n_1592);
 assign sub_1096_2_n_36 = ~(in1_128_8_ | ~n_1590);
 assign sub_1096_2_n_35 = ~(in1_128_20_ | ~n_1594);
 assign sub_1096_2_n_18 = ~sub_1096_2_n_17;
 assign sub_1096_2_n_13 = ~sub_1096_2_n_12;
 assign sub_1096_2_n_34 = ~(in1_128_6_ & ~n_1528);
 assign sub_1096_2_n_33 = ~(in1_128_20_ & ~n_1594);
 assign sub_1096_2_n_32 = ~(n_1496 | ~in1_128_14_);
 assign sub_1096_2_n_31 = ~(in1_128_22_ & ~n_1404);
 assign sub_1096_2_n_30 = ~(in1_128_4_ & ~n_1570);
 assign sub_1096_2_n_29 = ~(in1_128_12_ | ~n_1582);
 assign sub_1096_2_n_28 = ~(in1_128_15_ & ~n_1550);
 assign sub_1096_2_n_27 = ~(in1_128_17_ & ~n_1473);
 assign sub_1096_2_n_26 = ~(in1_128_10_ | ~n_1556);
 assign sub_1096_2_n_25 = ~(in1_128_3_ | ~n_1536);
 assign sub_1096_2_n_24 = ~(in1_128_14_ | ~n_1496);
 assign sub_1096_2_n_23 = ~(in1_128_4_ | ~n_1570);
 assign sub_1096_2_n_22 = ~(in1_128_3_ & ~n_1536);
 assign sub_1096_2_n_21 = ~(in1_128_7_ & ~n_1480);
 assign sub_1096_2_n_20 = ~(in1_128_9_ | ~n_1552);
 assign sub_1096_2_n_19 = ~(in1_128_15_ | ~n_1550);
 assign sub_1096_2_n_17 = ~(in1_128_1_ | ~n_1478);
 assign sub_1096_2_n_16 = ~(in1_128_21_ & ~n_1592);
 assign sub_1096_2_n_15 = ~(in1_128_19_ & ~n_1566);
 assign sub_1096_2_n_14 = ~(in1_128_18_ | ~n_1559);
 assign sub_1096_2_n_12 = ~(in1_128_1_ & ~n_1478);
 assign sub_1096_2_n_11 = ~(n_1544 & ~n_1574);
 assign sub_1096_2_n_10 = ~n_1587;
 assign sub_1096_2_n_9 = ~n_1544;
 assign sub_1096_2_n_8 = (sub_1096_2_n_131 & sub_1096_2_n_115);
 assign in1_130_22_ = ~(sub_1096_2_n_166 ^ sub_1096_2_n_86);
 assign sub_1096_2_n_6 = ~(sub_1096_2_n_70 & ~sub_1096_2_n_72);
 assign in1_130_15_ = (sub_1096_2_n_163 ^ sub_1096_2_n_69);
 assign sub_1096_2_n_4 = ~(sub_1096_2_n_8 | ~sub_1096_2_n_68);
 assign sub_1096_2_n_3 = ~(in1_128_2_ | ~n_1580);
 assign sub_1096_2_n_2 = ~(in1_128_13_ | ~n_1578);
 assign sub_1096_2_n_1 = ~(in1_128_16_ | ~n_1563);
 assign sub_1096_2_n_0 = ~(in1_128_5_ | ~n_1568);
 assign in1_133_23_ = ~(sub_1117_2_n_157 ^ sub_1117_2_n_74);
 assign sub_1117_2_n_157 = ~(sub_1117_2_n_10 & (sub_1117_2_n_152 | sub_1117_2_n_31));
 assign in1_133_22_ = ~(sub_1117_2_n_152 ^ sub_1117_2_n_70);
 assign in1_133_21_ = ~(sub_1117_2_n_151 ^ sub_1117_2_n_69);
 assign in1_133_19_ = ~(sub_1117_2_n_150 ^ sub_1117_2_n_57);
 assign in1_133_15_ = ~(sub_1117_2_n_146 ^ sub_1117_2_n_51);
 assign sub_1117_2_n_152 = ~(sub_1117_2_n_90 | (sub_1117_2_n_141 & sub_1117_2_n_67));
 assign sub_1117_2_n_151 = ~(sub_1117_2_n_4 & ~(sub_1117_2_n_141 & sub_1117_2_n_36));
 assign sub_1117_2_n_150 = ~(sub_1117_2_n_37 & (sub_1117_2_n_140 | sub_1117_2_n_43));
 assign in1_133_20_ = ~(sub_1117_2_n_141 ^ sub_1117_2_n_68);
 assign in1_133_18_ = ~(sub_1117_2_n_140 ^ sub_1117_2_n_50);
 assign in1_133_17_ = ~(sub_1117_2_n_139 ^ sub_1117_2_n_62);
 assign sub_1117_2_n_146 = ~(sub_1117_2_n_40 & (sub_1117_2_n_135 | sub_1117_2_n_18));
 assign in1_133_24_ = ~(sub_1117_2_n_136 ^ in1_131_23_);
 assign in1_133_14_ = ~(sub_1117_2_n_135 ^ sub_1117_2_n_56);
 assign in1_133_13_ = ~(sub_1117_2_n_134 ^ sub_1117_2_n_55);
 assign in1_133_11_ = ~(sub_1117_2_n_133 ^ sub_1117_2_n_52);
 assign sub_1117_2_n_141 = ~(sub_1117_2_n_104 & (sub_1117_2_n_129 | sub_1117_2_n_97));
 assign sub_1117_2_n_140 = ~(sub_1117_2_n_137 | sub_1117_2_n_89);
 assign sub_1117_2_n_139 = ~(sub_1117_2_n_7 & (sub_1117_2_n_129 | sub_1117_2_n_39));
 assign in1_133_16_ = ~(sub_1117_2_n_129 ^ sub_1117_2_n_60);
 assign sub_1117_2_n_137 = ~(sub_1117_2_n_129 | sub_1117_2_n_79);
 assign sub_1117_2_n_136 = ~(sub_1117_2_n_113 & (sub_1117_2_n_127 | sub_1117_2_n_99));
 assign sub_1117_2_n_135 = ~(sub_1117_2_n_96 | (sub_1117_2_n_126 & sub_1117_2_n_81));
 assign sub_1117_2_n_134 = ~(sub_1117_2_n_35 & ~(sub_1117_2_n_126 & sub_1117_2_n_14));
 assign sub_1117_2_n_133 = ~(sub_1117_2_n_44 & (sub_1117_2_n_125 | sub_1117_2_n_20));
 assign in1_133_12_ = ~(sub_1117_2_n_126 ^ sub_1117_2_n_54);
 assign in1_133_10_ = ~(sub_1117_2_n_125 ^ sub_1117_2_n_75);
 assign in1_133_9_ = ~(sub_1117_2_n_124 ^ sub_1117_2_n_73);
 assign sub_1117_2_n_129 = (sub_1117_2_n_127 & sub_1117_2_n_108);
 assign in1_133_7_ = ~(sub_1117_2_n_122 ^ sub_1117_2_n_59);
 assign sub_1117_2_n_127 = ~(sub_1117_2_n_0 & sub_1117_2_n_95);
 assign sub_1117_2_n_126 = (sub_1117_2_n_0 | sub_1117_2_n_103);
 assign sub_1117_2_n_125 = ~(sub_1117_2_n_88 | (sub_1117_2_n_119 & sub_1117_2_n_65));
 assign sub_1117_2_n_124 = ~(sub_1117_2_n_29 & ~(sub_1117_2_n_119 & sub_1117_2_n_12));
 assign in1_133_8_ = ~(sub_1117_2_n_119 ^ sub_1117_2_n_53);
 assign sub_1117_2_n_122 = ~(sub_1117_2_n_34 & (sub_1117_2_n_118 | sub_1117_2_n_38));
 assign in1_133_6_ = ~(sub_1117_2_n_118 ^ sub_1117_2_n_61);
 assign in1_133_5_ = ~(sub_1117_2_n_117 ^ sub_1117_2_n_71);
 assign sub_1117_2_n_119 = ~(sub_1117_2_n_102 & ~(sub_1117_2_n_114 & sub_1117_2_n_83));
 assign sub_1117_2_n_118 = ~(sub_1117_2_n_114 | sub_1117_2_n_91);
 assign sub_1117_2_n_117 = ~(sub_1117_2_n_41 & (sub_1117_2_n_109 | sub_1117_2_n_5));
 assign in1_133_4_ = ~(sub_1117_2_n_109 ^ sub_1117_2_n_72);
 assign in1_133_3_ = ~(sub_1117_2_n_111 ^ sub_1117_2_n_58);
 assign sub_1117_2_n_114 = ~(sub_1117_2_n_109 | sub_1117_2_n_77);
 assign sub_1117_2_n_113 = ~sub_1117_2_n_112;
 assign sub_1117_2_n_112 = ~(sub_1117_2_n_105 & (sub_1117_2_n_100 & (sub_1117_2_n_108 | sub_1117_2_n_99)));
 assign sub_1117_2_n_111 = ~(sub_1117_2_n_33 | (sub_1117_2_n_107 & sub_1117_2_n_9));
 assign in1_133_2_ = ~(sub_1117_2_n_107 ^ sub_1117_2_n_76);
 assign sub_1117_2_n_109 = ~(sub_1117_2_n_85 | (sub_1117_2_n_107 & sub_1117_2_n_64));
 assign sub_1117_2_n_108 = ~(sub_1117_2_n_101 | (sub_1117_2_n_103 & sub_1117_2_n_95));
 assign sub_1117_2_n_107 = ((sub_1117_2_n_3 & in1_131_0_) | ((in1_131_0_ & sub_1117_2_n_2) | (sub_1117_2_n_2
    & sub_1117_2_n_3)));
 assign in1_133_1_ = (in1_131_0_ ^ (sub_1117_2_n_2 ^ sub_1117_2_n_3));
 assign sub_1117_2_n_105 = ~(sub_1117_2_n_98 & ~sub_1117_2_n_104);
 assign sub_1117_2_n_104 = ~(sub_1117_2_n_93 | (sub_1117_2_n_89 & sub_1117_2_n_80));
 assign sub_1117_2_n_103 = ~(sub_1117_2_n_86 & ~(sub_1117_2_n_88 & sub_1117_2_n_66));
 assign sub_1117_2_n_102 = ~(sub_1117_2_n_78 | (sub_1117_2_n_45 | (sub_1117_2_n_91 & sub_1117_2_n_83)));
 assign sub_1117_2_n_101 = ~(sub_1117_2_n_92 & ~(sub_1117_2_n_96 & sub_1117_2_n_84));
 assign sub_1117_2_n_100 = ~(sub_1117_2_n_87 | (sub_1117_2_n_90 & sub_1117_2_n_82));
 assign sub_1117_2_n_99 = ~(sub_1117_2_n_98 & ~sub_1117_2_n_97);
 assign sub_1117_2_n_94 = ~(sub_1117_2_n_65 & sub_1117_2_n_66);
 assign sub_1117_2_n_93 = ~(sub_1117_2_n_24 & (sub_1117_2_n_37 | sub_1117_2_n_19));
 assign sub_1117_2_n_92 = ~(sub_1117_2_n_23 | ~(sub_1117_2_n_40 | sub_1117_2_n_30));
 assign sub_1117_2_n_98 = (sub_1117_2_n_67 & sub_1117_2_n_82);
 assign sub_1117_2_n_97 = ~(sub_1117_2_n_80 & ~sub_1117_2_n_79);
 assign sub_1117_2_n_96 = ~(sub_1117_2_n_48 & (sub_1117_2_n_35 | sub_1117_2_n_42));
 assign sub_1117_2_n_95 = (sub_1117_2_n_81 & sub_1117_2_n_84);
 assign sub_1117_2_n_87 = ~(sub_1117_2_n_25 & (sub_1117_2_n_10 | sub_1117_2_n_15));
 assign sub_1117_2_n_86 = ~(sub_1117_2_n_47 | ~(sub_1117_2_n_44 | sub_1117_2_n_6));
 assign sub_1117_2_n_85 = ~(sub_1117_2_n_46 & (sub_1117_2_n_32 | sub_1117_2_n_13));
 assign sub_1117_2_n_91 = ~(sub_1117_2_n_49 & (sub_1117_2_n_41 | sub_1117_2_n_11));
 assign sub_1117_2_n_90 = ~(sub_1117_2_n_21 & (sub_1117_2_n_4 | sub_1117_2_n_16));
 assign sub_1117_2_n_89 = ~(sub_1117_2_n_22 & (sub_1117_2_n_7 | sub_1117_2_n_17));
 assign sub_1117_2_n_88 = ~(sub_1117_2_n_26 & (sub_1117_2_n_29 | sub_1117_2_n_28));
 assign sub_1117_2_n_78 = ~(sub_1117_2_n_34 | sub_1117_2_n_27);
 assign sub_1117_2_n_77 = (sub_1117_2_n_5 | sub_1117_2_n_11);
 assign sub_1117_2_n_76 = ~(sub_1117_2_n_32 & sub_1117_2_n_9);
 assign sub_1117_2_n_75 = ~(sub_1117_2_n_20 | ~sub_1117_2_n_44);
 assign sub_1117_2_n_84 = ~(sub_1117_2_n_18 | sub_1117_2_n_30);
 assign sub_1117_2_n_83 = ~(sub_1117_2_n_38 | sub_1117_2_n_27);
 assign sub_1117_2_n_74 = ~(sub_1117_2_n_25 & ~sub_1117_2_n_15);
 assign sub_1117_2_n_73 = ~(sub_1117_2_n_26 & ~sub_1117_2_n_28);
 assign sub_1117_2_n_72 = ~(sub_1117_2_n_5 | ~sub_1117_2_n_41);
 assign sub_1117_2_n_82 = ~(sub_1117_2_n_31 | sub_1117_2_n_15);
 assign sub_1117_2_n_71 = ~(sub_1117_2_n_49 & ~sub_1117_2_n_11);
 assign sub_1117_2_n_70 = ~(sub_1117_2_n_31 | ~sub_1117_2_n_10);
 assign sub_1117_2_n_69 = ~(sub_1117_2_n_21 & ~sub_1117_2_n_16);
 assign sub_1117_2_n_81 = ~(sub_1117_2_n_42 | ~sub_1117_2_n_14);
 assign sub_1117_2_n_80 = ~(sub_1117_2_n_43 | sub_1117_2_n_19);
 assign sub_1117_2_n_79 = (sub_1117_2_n_39 | sub_1117_2_n_17);
 assign sub_1117_2_n_68 = ~(sub_1117_2_n_4 & sub_1117_2_n_36);
 assign sub_1117_2_n_64 = ~(sub_1117_2_n_8 | sub_1117_2_n_13);
 assign in1_133_0_ = ~(sub_1117_2_n_3 & ~(sub_1117_2_n_1 & n_1531));
 assign sub_1117_2_n_62 = ~(sub_1117_2_n_22 & ~sub_1117_2_n_17);
 assign sub_1117_2_n_61 = ~(sub_1117_2_n_38 | ~sub_1117_2_n_34);
 assign sub_1117_2_n_60 = ~(sub_1117_2_n_39 | ~sub_1117_2_n_7);
 assign sub_1117_2_n_59 = (sub_1117_2_n_45 | sub_1117_2_n_27);
 assign sub_1117_2_n_67 = ~(sub_1117_2_n_16 | ~sub_1117_2_n_36);
 assign sub_1117_2_n_58 = ~(sub_1117_2_n_13 | ~sub_1117_2_n_46);
 assign sub_1117_2_n_66 = ~(sub_1117_2_n_20 | sub_1117_2_n_6);
 assign sub_1117_2_n_57 = ~(sub_1117_2_n_24 & ~sub_1117_2_n_19);
 assign sub_1117_2_n_56 = ~(sub_1117_2_n_18 | ~sub_1117_2_n_40);
 assign sub_1117_2_n_55 = ~(sub_1117_2_n_48 & ~sub_1117_2_n_42);
 assign sub_1117_2_n_54 = ~(sub_1117_2_n_35 & sub_1117_2_n_14);
 assign sub_1117_2_n_53 = ~(sub_1117_2_n_29 & sub_1117_2_n_12);
 assign sub_1117_2_n_52 = (sub_1117_2_n_47 | sub_1117_2_n_6);
 assign sub_1117_2_n_51 = (sub_1117_2_n_23 | sub_1117_2_n_30);
 assign sub_1117_2_n_65 = ~(sub_1117_2_n_28 | ~sub_1117_2_n_12);
 assign sub_1117_2_n_50 = ~(sub_1117_2_n_43 | ~sub_1117_2_n_37);
 assign sub_1117_2_n_33 = ~sub_1117_2_n_32;
 assign sub_1117_2_n_49 = ~(in1_131_4_ & ~n_1570);
 assign sub_1117_2_n_48 = ~(in1_131_12_ & ~n_1582);
 assign sub_1117_2_n_47 = ~(n_1556 | ~in1_131_10_);
 assign sub_1117_2_n_46 = ~(in1_131_2_ & ~n_1580);
 assign sub_1117_2_n_45 = ~(n_1528 | ~in1_131_6_);
 assign sub_1117_2_n_44 = ~(in1_131_9_ & ~n_1552);
 assign sub_1117_2_n_43 = ~(in1_131_17_ | ~n_1473);
 assign sub_1117_2_n_42 = ~(in1_131_12_ | ~n_1582);
 assign sub_1117_2_n_41 = ~(in1_131_3_ & ~n_1536);
 assign sub_1117_2_n_40 = ~(in1_131_13_ & ~n_1578);
 assign sub_1117_2_n_39 = ~(in1_131_15_ | ~n_1550);
 assign sub_1117_2_n_38 = ~(in1_131_5_ | ~n_1568);
 assign sub_1117_2_n_37 = ~(in1_131_17_ & ~n_1473);
 assign sub_1117_2_n_36 = ~(n_1566 & ~in1_131_19_);
 assign sub_1117_2_n_35 = ~(in1_131_11_ & ~n_1596);
 assign sub_1117_2_n_34 = ~(in1_131_5_ & ~n_1568);
 assign sub_1117_2_n_32 = ~(in1_131_1_ & ~n_1478);
 assign sub_1117_2_n_31 = ~(in1_131_21_ | ~n_1592);
 assign sub_1117_2_n_30 = ~(in1_131_14_ | ~n_1496);
 assign sub_1117_2_n_29 = ~(in1_131_7_ & ~n_1480);
 assign sub_1117_2_n_28 = ~(in1_131_8_ | ~n_1590);
 assign sub_1117_2_n_27 = ~(in1_131_6_ | ~n_1528);
 assign sub_1117_2_n_9 = ~sub_1117_2_n_8;
 assign sub_1117_2_n_26 = ~(in1_131_8_ & ~n_1590);
 assign sub_1117_2_n_25 = ~(in1_131_22_ & ~n_1404);
 assign sub_1117_2_n_24 = ~(in1_131_18_ & ~n_1559);
 assign sub_1117_2_n_23 = ~(n_1496 | ~in1_131_14_);
 assign sub_1117_2_n_22 = ~(in1_131_16_ & ~n_1563);
 assign sub_1117_2_n_21 = ~(in1_131_20_ & ~n_1594);
 assign sub_1117_2_n_20 = ~(in1_131_9_ | ~n_1552);
 assign sub_1117_2_n_19 = ~(in1_131_18_ | ~n_1559);
 assign sub_1117_2_n_18 = ~(in1_131_13_ | ~n_1578);
 assign sub_1117_2_n_17 = ~(in1_131_16_ | ~n_1563);
 assign sub_1117_2_n_16 = ~(in1_131_20_ | ~n_1594);
 assign sub_1117_2_n_15 = ~(in1_131_22_ | ~n_1404);
 assign sub_1117_2_n_14 = ~(n_1596 & ~in1_131_11_);
 assign sub_1117_2_n_13 = ~(in1_131_2_ | ~n_1580);
 assign sub_1117_2_n_12 = ~(n_1480 & ~in1_131_7_);
 assign sub_1117_2_n_11 = ~(in1_131_4_ | ~n_1570);
 assign sub_1117_2_n_10 = ~(in1_131_21_ & ~n_1592);
 assign sub_1117_2_n_8 = ~(in1_131_1_ | ~n_1478);
 assign sub_1117_2_n_7 = ~(in1_131_15_ & ~n_1550);
 assign sub_1117_2_n_6 = ~(in1_131_10_ | ~n_1556);
 assign sub_1117_2_n_5 = ~(in1_131_3_ | ~n_1536);
 assign sub_1117_2_n_4 = ~(in1_131_19_ & ~n_1566);
 assign sub_1117_2_n_3 = ~(n_1544 & ~n_1531);
 assign sub_1117_2_n_2 = ~n_1587;
 assign sub_1117_2_n_1 = ~n_1544;
 assign sub_1117_2_n_0 = ~(sub_1117_2_n_94 | ~sub_1117_2_n_119);
 assign in1_136_23_ = ~(sub_1138_2_n_151 ^ sub_1138_2_n_73);
 assign sub_1138_2_n_151 = ~(sub_1138_2_n_6 & (sub_1138_2_n_146 | sub_1138_2_n_30));
 assign in1_136_22_ = ~(sub_1138_2_n_146 ^ sub_1138_2_n_70);
 assign in1_136_21_ = ~(sub_1138_2_n_145 ^ sub_1138_2_n_69);
 assign in1_136_19_ = ~(sub_1138_2_n_144 ^ sub_1138_2_n_66);
 assign in1_136_15_ = ~(sub_1138_2_n_143 ^ sub_1138_2_n_56);
 assign sub_1138_2_n_146 = ~(sub_1138_2_n_84 | (sub_1138_2_n_135 & sub_1138_2_n_77));
 assign sub_1138_2_n_145 = ~(sub_1138_2_n_5 & ~(sub_1138_2_n_135 & sub_1138_2_n_39));
 assign sub_1138_2_n_144 = ~(sub_1138_2_n_18 & (sub_1138_2_n_134 | sub_1138_2_n_34));
 assign sub_1138_2_n_143 = ~(sub_1138_2_n_42 & (sub_1138_2_n_132 | sub_1138_2_n_26));
 assign in1_136_20_ = ~(sub_1138_2_n_135 ^ sub_1138_2_n_68);
 assign in1_136_18_ = ~(sub_1138_2_n_134 ^ sub_1138_2_n_57);
 assign in1_136_17_ = ~(sub_1138_2_n_133 ^ sub_1138_2_n_60);
 assign in1_136_14_ = ~(sub_1138_2_n_132 ^ sub_1138_2_n_54);
 assign in1_136_13_ = ~(sub_1138_2_n_131 ^ sub_1138_2_n_53);
 assign in1_136_11_ = ~(sub_1138_2_n_130 ^ sub_1138_2_n_59);
 assign in1_136_24_ = ~(sub_1138_2_n_125 ^ in1_134_23_);
 assign sub_1138_2_n_135 = ~(sub_1138_2_n_96 & (sub_1138_2_n_123 | sub_1138_2_n_90));
 assign sub_1138_2_n_134 = ~(sub_1138_2_n_83 | ~(sub_1138_2_n_123 | sub_1138_2_n_63));
 assign sub_1138_2_n_133 = ~(sub_1138_2_n_19 & (sub_1138_2_n_123 | sub_1138_2_n_8));
 assign sub_1138_2_n_132 = ~(sub_1138_2_n_87 | (sub_1138_2_n_122 & sub_1138_2_n_78));
 assign sub_1138_2_n_131 = ~(sub_1138_2_n_38 & ~(sub_1138_2_n_122 & sub_1138_2_n_31));
 assign sub_1138_2_n_130 = ~(sub_1138_2_n_33 & (sub_1138_2_n_121 | sub_1138_2_n_9));
 assign in1_136_16_ = ~(sub_1138_2_n_123 ^ sub_1138_2_n_75);
 assign in1_136_12_ = ~(sub_1138_2_n_122 ^ sub_1138_2_n_50);
 assign in1_136_10_ = ~(sub_1138_2_n_121 ^ sub_1138_2_n_51);
 assign in1_136_9_ = ~(sub_1138_2_n_120 ^ sub_1138_2_n_72);
 assign sub_1138_2_n_125 = ~(sub_1138_2_n_103 & ((sub_1138_2_n_104 | sub_1138_2_n_93) & (sub_1138_2_n_117
    | sub_1138_2_n_93)));
 assign in1_136_7_ = ~(sub_1138_2_n_118 ^ sub_1138_2_n_55);
 assign sub_1138_2_n_123 = (sub_1138_2_n_117 & sub_1138_2_n_104);
 assign sub_1138_2_n_122 = ~(sub_1138_2_n_99 & (sub_1138_2_n_113 | sub_1138_2_n_89));
 assign sub_1138_2_n_121 = ~(sub_1138_2_n_86 | (sub_1138_2_n_114 & sub_1138_2_n_64));
 assign sub_1138_2_n_120 = ~(sub_1138_2_n_10 & (sub_1138_2_n_113 | sub_1138_2_n_36));
 assign in1_136_8_ = ~(sub_1138_2_n_114 ^ sub_1138_2_n_74);
 assign sub_1138_2_n_118 = ~(sub_1138_2_n_35 & (sub_1138_2_n_112 | sub_1138_2_n_40));
 assign sub_1138_2_n_117 = ~(sub_1138_2_n_91 & (sub_1138_2_n_114 & ~sub_1138_2_n_89));
 assign in1_136_6_ = ~(sub_1138_2_n_112 ^ sub_1138_2_n_71);
 assign in1_136_5_ = ~(sub_1138_2_n_111 ^ sub_1138_2_n_52);
 assign sub_1138_2_n_113 = ~sub_1138_2_n_114;
 assign sub_1138_2_n_114 = ~(sub_1138_2_n_98 & ~(sub_1138_2_n_108 & sub_1138_2_n_82));
 assign sub_1138_2_n_112 = ~(sub_1138_2_n_108 | sub_1138_2_n_85);
 assign sub_1138_2_n_111 = ~(sub_1138_2_n_11 & (sub_1138_2_n_105 | sub_1138_2_n_14));
 assign in1_136_4_ = ~(sub_1138_2_n_105 ^ sub_1138_2_n_49);
 assign in1_136_3_ = ~(sub_1138_2_n_107 ^ sub_1138_2_n_58);
 assign sub_1138_2_n_108 = ~(sub_1138_2_n_14 | (sub_1138_2_n_12 | sub_1138_2_n_105));
 assign sub_1138_2_n_107 = ~(sub_1138_2_n_3 | (sub_1138_2_n_102 & sub_1138_2_n_7));
 assign in1_136_2_ = ~(sub_1138_2_n_102 ^ sub_1138_2_n_67);
 assign sub_1138_2_n_105 = ~(sub_1138_2_n_48 | ((sub_1138_2_n_102 & sub_1138_2_n_62) | (sub_1138_2_n_3
    & sub_1138_2_n_16)));
 assign sub_1138_2_n_104 = ~(sub_1138_2_n_100 | sub_1138_2_n_97);
 assign sub_1138_2_n_103 = ~(sub_1138_2_n_95 | ~(sub_1138_2_n_96 | sub_1138_2_n_88));
 assign sub_1138_2_n_102 = ((sub_1138_2_n_2 & in1_134_0_) | ((in1_134_0_ & sub_1138_2_n_1) | (sub_1138_2_n_1
    & sub_1138_2_n_2)));
 assign in1_136_1_ = (in1_134_0_ ^ (sub_1138_2_n_1 ^ sub_1138_2_n_2));
 assign sub_1138_2_n_100 = ~(sub_1138_2_n_99 | ~sub_1138_2_n_91);
 assign sub_1138_2_n_99 = ~(sub_1138_2_n_46 | ((sub_1138_2_n_86 & sub_1138_2_n_65) | (sub_1138_2_n_32
    & sub_1138_2_n_15)));
 assign sub_1138_2_n_98 = ~(sub_1138_2_n_76 | (sub_1138_2_n_25 | (sub_1138_2_n_85 & sub_1138_2_n_82)));
 assign sub_1138_2_n_97 = ~(sub_1138_2_n_23 & (sub_1138_2_n_94 & (sub_1138_2_n_42 | sub_1138_2_n_13)));
 assign sub_1138_2_n_96 = ~(sub_1138_2_n_47 | ((sub_1138_2_n_83 & sub_1138_2_n_79) | (sub_1138_2_n_17
    & sub_1138_2_n_4)));
 assign sub_1138_2_n_95 = ~(sub_1138_2_n_22 & (sub_1138_2_n_92 & (sub_1138_2_n_6 | sub_1138_2_n_41)));
 assign sub_1138_2_n_94 = ~(sub_1138_2_n_87 & sub_1138_2_n_81);
 assign sub_1138_2_n_93 = (sub_1138_2_n_90 | sub_1138_2_n_88);
 assign sub_1138_2_n_92 = ~(sub_1138_2_n_84 & sub_1138_2_n_80);
 assign sub_1138_2_n_91 = (sub_1138_2_n_78 & sub_1138_2_n_81);
 assign sub_1138_2_n_90 = ~(sub_1138_2_n_79 & ~sub_1138_2_n_63);
 assign sub_1138_2_n_89 = ~(sub_1138_2_n_64 & sub_1138_2_n_65);
 assign sub_1138_2_n_88 = ~(sub_1138_2_n_77 & sub_1138_2_n_80);
 assign sub_1138_2_n_87 = ~(sub_1138_2_n_45 & (sub_1138_2_n_38 | sub_1138_2_n_20));
 assign sub_1138_2_n_86 = ~(sub_1138_2_n_44 & (sub_1138_2_n_10 | sub_1138_2_n_29));
 assign sub_1138_2_n_85 = ~(sub_1138_2_n_21 & (sub_1138_2_n_11 | sub_1138_2_n_12));
 assign sub_1138_2_n_84 = ~(sub_1138_2_n_24 & (sub_1138_2_n_5 | sub_1138_2_n_27));
 assign sub_1138_2_n_83 = ~(sub_1138_2_n_43 & (sub_1138_2_n_19 | sub_1138_2_n_28));
 assign sub_1138_2_n_76 = ~(sub_1138_2_n_35 | sub_1138_2_n_37);
 assign sub_1138_2_n_75 = ~(sub_1138_2_n_8 | ~sub_1138_2_n_19);
 assign sub_1138_2_n_74 = ~(sub_1138_2_n_10 & ~sub_1138_2_n_36);
 assign sub_1138_2_n_73 = ~(sub_1138_2_n_22 & ~sub_1138_2_n_41);
 assign sub_1138_2_n_82 = ~(sub_1138_2_n_40 | sub_1138_2_n_37);
 assign sub_1138_2_n_72 = ~(sub_1138_2_n_44 & ~sub_1138_2_n_29);
 assign sub_1138_2_n_81 = ~(sub_1138_2_n_26 | sub_1138_2_n_13);
 assign sub_1138_2_n_71 = ~(sub_1138_2_n_40 | ~sub_1138_2_n_35);
 assign sub_1138_2_n_80 = ~(sub_1138_2_n_30 | sub_1138_2_n_41);
 assign sub_1138_2_n_70 = ~(sub_1138_2_n_30 | ~sub_1138_2_n_6);
 assign sub_1138_2_n_69 = ~(sub_1138_2_n_24 & ~sub_1138_2_n_27);
 assign sub_1138_2_n_79 = ~(sub_1138_2_n_34 | ~sub_1138_2_n_4);
 assign sub_1138_2_n_78 = ~(sub_1138_2_n_20 | ~sub_1138_2_n_31);
 assign sub_1138_2_n_68 = ~(sub_1138_2_n_5 & sub_1138_2_n_39);
 assign sub_1138_2_n_67 = ~(sub_1138_2_n_7 & ~sub_1138_2_n_3);
 assign sub_1138_2_n_66 = ~(sub_1138_2_n_4 & ~sub_1138_2_n_47);
 assign sub_1138_2_n_77 = ~(sub_1138_2_n_27 | ~sub_1138_2_n_39);
 assign sub_1138_2_n_62 = (sub_1138_2_n_7 & sub_1138_2_n_16);
 assign in1_136_0_ = ~(sub_1138_2_n_2 & ~(sub_1138_2_n_0 & n_1554));
 assign sub_1138_2_n_60 = ~(sub_1138_2_n_43 & ~sub_1138_2_n_28);
 assign sub_1138_2_n_59 = ~(sub_1138_2_n_15 & ~sub_1138_2_n_46);
 assign sub_1138_2_n_65 = ~(sub_1138_2_n_9 | ~sub_1138_2_n_15);
 assign sub_1138_2_n_64 = ~(sub_1138_2_n_36 | sub_1138_2_n_29);
 assign sub_1138_2_n_58 = ~(sub_1138_2_n_48 | ~sub_1138_2_n_16);
 assign sub_1138_2_n_57 = ~(sub_1138_2_n_17 | sub_1138_2_n_34);
 assign sub_1138_2_n_56 = ~(sub_1138_2_n_23 & ~sub_1138_2_n_13);
 assign sub_1138_2_n_55 = (sub_1138_2_n_25 | sub_1138_2_n_37);
 assign sub_1138_2_n_54 = ~(sub_1138_2_n_26 | ~sub_1138_2_n_42);
 assign sub_1138_2_n_53 = ~(sub_1138_2_n_45 & ~sub_1138_2_n_20);
 assign sub_1138_2_n_52 = ~(sub_1138_2_n_21 & ~sub_1138_2_n_12);
 assign sub_1138_2_n_63 = (sub_1138_2_n_8 | sub_1138_2_n_28);
 assign sub_1138_2_n_51 = ~(sub_1138_2_n_32 | sub_1138_2_n_9);
 assign sub_1138_2_n_50 = ~(sub_1138_2_n_38 & sub_1138_2_n_31);
 assign sub_1138_2_n_49 = ~(sub_1138_2_n_14 | ~sub_1138_2_n_11);
 assign sub_1138_2_n_33 = ~sub_1138_2_n_32;
 assign sub_1138_2_n_48 = ~(n_1580 | ~in1_134_2_);
 assign sub_1138_2_n_47 = ~(n_1559 | ~in1_134_18_);
 assign sub_1138_2_n_46 = ~(n_1556 | ~in1_134_10_);
 assign sub_1138_2_n_45 = ~(in1_134_12_ & ~n_1582);
 assign sub_1138_2_n_44 = ~(in1_134_8_ & ~n_1590);
 assign sub_1138_2_n_43 = ~(in1_134_16_ & ~n_1563);
 assign sub_1138_2_n_42 = ~(in1_134_13_ & ~n_1578);
 assign sub_1138_2_n_41 = ~(in1_134_22_ | ~n_1404);
 assign sub_1138_2_n_40 = ~(in1_134_5_ | ~n_1568);
 assign sub_1138_2_n_39 = ~(n_1566 & ~in1_134_19_);
 assign sub_1138_2_n_38 = ~(in1_134_11_ & ~n_1596);
 assign sub_1138_2_n_37 = ~(in1_134_6_ | ~n_1528);
 assign sub_1138_2_n_36 = ~(in1_134_7_ | ~n_1480);
 assign sub_1138_2_n_35 = ~(in1_134_5_ & ~n_1568);
 assign sub_1138_2_n_34 = ~(in1_134_17_ | ~n_1473);
 assign sub_1138_2_n_32 = ~(n_1552 | ~in1_134_9_);
 assign sub_1138_2_n_31 = ~(n_1596 & ~in1_134_11_);
 assign sub_1138_2_n_30 = ~(in1_134_21_ | ~n_1592);
 assign sub_1138_2_n_29 = ~(in1_134_8_ | ~n_1590);
 assign sub_1138_2_n_28 = ~(in1_134_16_ | ~n_1563);
 assign sub_1138_2_n_27 = ~(in1_134_20_ | ~n_1594);
 assign sub_1138_2_n_26 = ~(in1_134_13_ | ~n_1578);
 assign sub_1138_2_n_18 = ~sub_1138_2_n_17;
 assign sub_1138_2_n_25 = ~(n_1528 | ~in1_134_6_);
 assign sub_1138_2_n_24 = ~(in1_134_20_ & ~n_1594);
 assign sub_1138_2_n_23 = ~(in1_134_14_ & ~n_1496);
 assign sub_1138_2_n_22 = ~(in1_134_22_ & ~n_1404);
 assign sub_1138_2_n_21 = ~(in1_134_4_ & ~n_1570);
 assign sub_1138_2_n_20 = ~(in1_134_12_ | ~n_1582);
 assign sub_1138_2_n_19 = ~(in1_134_15_ & ~n_1550);
 assign sub_1138_2_n_17 = ~(n_1473 | ~in1_134_17_);
 assign sub_1138_2_n_16 = ~(n_1580 & ~in1_134_2_);
 assign sub_1138_2_n_15 = ~(n_1556 & ~in1_134_10_);
 assign sub_1138_2_n_14 = ~(in1_134_3_ | ~n_1536);
 assign sub_1138_2_n_13 = ~(in1_134_14_ | ~n_1496);
 assign sub_1138_2_n_12 = ~(in1_134_4_ | ~n_1570);
 assign sub_1138_2_n_11 = ~(in1_134_3_ & ~n_1536);
 assign sub_1138_2_n_10 = ~(in1_134_7_ & ~n_1480);
 assign sub_1138_2_n_9 = ~(in1_134_9_ | ~n_1552);
 assign sub_1138_2_n_8 = ~(in1_134_15_ | ~n_1550);
 assign sub_1138_2_n_7 = ~(n_1478 & ~in1_134_1_);
 assign sub_1138_2_n_6 = ~(in1_134_21_ & ~n_1592);
 assign sub_1138_2_n_5 = ~(in1_134_19_ & ~n_1566);
 assign sub_1138_2_n_4 = ~(n_1559 & ~in1_134_18_);
 assign sub_1138_2_n_3 = ~(n_1478 | ~in1_134_1_);
 assign sub_1138_2_n_2 = ~(n_1544 & ~n_1554);
 assign sub_1138_2_n_1 = ~n_1587;
 assign sub_1138_2_n_0 = ~n_1544;
 assign in1_139_23_ = ~(sub_1159_2_n_147 ^ sub_1159_2_n_72);
 assign sub_1159_2_n_147 = ~(sub_1159_2_n_8 & (sub_1159_2_n_142 | sub_1159_2_n_29));
 assign in1_139_22_ = ~(sub_1159_2_n_142 ^ sub_1159_2_n_68);
 assign in1_139_21_ = ~(sub_1159_2_n_141 ^ sub_1159_2_n_67);
 assign in1_139_19_ = ~(sub_1159_2_n_140 ^ sub_1159_2_n_74);
 assign in1_139_15_ = ~(sub_1159_2_n_136 ^ sub_1159_2_n_49);
 assign sub_1159_2_n_142 = ~(sub_1159_2_n_81 | (sub_1159_2_n_131 & sub_1159_2_n_63));
 assign sub_1159_2_n_141 = ~(sub_1159_2_n_3 & ~(sub_1159_2_n_131 & sub_1159_2_n_33));
 assign sub_1159_2_n_140 = ~(sub_1159_2_n_35 & (sub_1159_2_n_130 | sub_1159_2_n_41));
 assign in1_139_20_ = ~(sub_1159_2_n_131 ^ sub_1159_2_n_66);
 assign in1_139_18_ = ~(sub_1159_2_n_130 ^ sub_1159_2_n_56);
 assign in1_139_17_ = ~(sub_1159_2_n_129 ^ sub_1159_2_n_48);
 assign sub_1159_2_n_136 = ~(sub_1159_2_n_38 & (sub_1159_2_n_126 | sub_1159_2_n_16));
 assign in1_139_24_ = ~(sub_1159_2_n_127 ^ in1_137_23_);
 assign in1_139_14_ = ~(sub_1159_2_n_126 ^ sub_1159_2_n_54);
 assign in1_139_13_ = ~(sub_1159_2_n_125 ^ sub_1159_2_n_53);
 assign in1_139_11_ = ~(sub_1159_2_n_124 ^ sub_1159_2_n_50);
 assign sub_1159_2_n_131 = ~(sub_1159_2_n_96 & (sub_1159_2_n_120 | sub_1159_2_n_88));
 assign sub_1159_2_n_130 = ~(sub_1159_2_n_82 | ~(sub_1159_2_n_120 | sub_1159_2_n_80));
 assign sub_1159_2_n_129 = ~(sub_1159_2_n_6 & (sub_1159_2_n_120 | sub_1159_2_n_37));
 assign in1_139_16_ = ~(sub_1159_2_n_120 ^ sub_1159_2_n_58);
 assign sub_1159_2_n_127 = ~(sub_1159_2_n_99 & ((sub_1159_2_n_100 | sub_1159_2_n_92) & (sub_1159_2_n_118
    | sub_1159_2_n_92)));
 assign sub_1159_2_n_126 = ~(sub_1159_2_n_83 | (sub_1159_2_n_117 & sub_1159_2_n_76));
 assign sub_1159_2_n_125 = ~(sub_1159_2_n_32 & ~(sub_1159_2_n_117 & sub_1159_2_n_12));
 assign sub_1159_2_n_124 = ~(sub_1159_2_n_42 & (sub_1159_2_n_116 | sub_1159_2_n_18));
 assign in1_139_12_ = ~(sub_1159_2_n_117 ^ sub_1159_2_n_52);
 assign in1_139_10_ = ~(sub_1159_2_n_116 ^ sub_1159_2_n_65);
 assign in1_139_9_ = ~(sub_1159_2_n_115 ^ sub_1159_2_n_71);
 assign sub_1159_2_n_120 = (sub_1159_2_n_118 & sub_1159_2_n_100);
 assign in1_139_7_ = ~(sub_1159_2_n_113 ^ sub_1159_2_n_57);
 assign sub_1159_2_n_118 = ~(sub_1159_2_n_112 & sub_1159_2_n_90);
 assign sub_1159_2_n_117 = (sub_1159_2_n_112 | sub_1159_2_n_95);
 assign sub_1159_2_n_116 = ~(sub_1159_2_n_84 | (sub_1159_2_n_109 & sub_1159_2_n_62));
 assign sub_1159_2_n_115 = ~(sub_1159_2_n_27 & ~(sub_1159_2_n_109 & sub_1159_2_n_10));
 assign in1_139_8_ = ~(sub_1159_2_n_109 ^ sub_1159_2_n_51);
 assign sub_1159_2_n_113 = ~(sub_1159_2_n_31 & (sub_1159_2_n_108 | sub_1159_2_n_36));
 assign sub_1159_2_n_112 = (sub_1159_2_n_62 & (sub_1159_2_n_64 & sub_1159_2_n_109));
 assign in1_139_6_ = ~(sub_1159_2_n_108 ^ sub_1159_2_n_59);
 assign in1_139_5_ = ~(sub_1159_2_n_107 ^ sub_1159_2_n_69);
 assign sub_1159_2_n_109 = ~(sub_1159_2_n_87 & ((sub_1159_2_n_85 | sub_1159_2_n_78) & (sub_1159_2_n_104
    | sub_1159_2_n_78)));
 assign sub_1159_2_n_108 = (sub_1159_2_n_104 & sub_1159_2_n_85);
 assign sub_1159_2_n_107 = ~(sub_1159_2_n_39 & (sub_1159_2_n_101 | sub_1159_2_n_4));
 assign in1_139_4_ = ~(sub_1159_2_n_101 ^ sub_1159_2_n_70);
 assign in1_139_3_ = ~(sub_1159_2_n_103 ^ sub_1159_2_n_55);
 assign sub_1159_2_n_104 = (sub_1159_2_n_4 | (sub_1159_2_n_9 | sub_1159_2_n_101));
 assign sub_1159_2_n_103 = ~(sub_1159_2_n_30 | (sub_1159_2_n_98 & sub_1159_2_n_7));
 assign in1_139_2_ = ~(sub_1159_2_n_98 ^ sub_1159_2_n_73);
 assign sub_1159_2_n_101 = ~(sub_1159_2_n_44 | ((sub_1159_2_n_98 & sub_1159_2_n_61) | (sub_1159_2_n_30
    & sub_1159_2_n_11)));
 assign sub_1159_2_n_100 = ~(sub_1159_2_n_86 | ((sub_1159_2_n_95 & sub_1159_2_n_90) | (sub_1159_2_n_83
    & sub_1159_2_n_79)));
 assign sub_1159_2_n_99 = ~(sub_1159_2_n_94 | ~(sub_1159_2_n_96 | sub_1159_2_n_89));
 assign sub_1159_2_n_98 = ((sub_1159_2_n_2 & in1_137_0_) | ((in1_137_0_ & sub_1159_2_n_1) | (sub_1159_2_n_1
    & sub_1159_2_n_2)));
 assign in1_139_1_ = (in1_137_0_ ^ (sub_1159_2_n_1 ^ sub_1159_2_n_2));
 assign sub_1159_2_n_96 = ~(sub_1159_2_n_22 | ((sub_1159_2_n_82 & sub_1159_2_n_75) | (sub_1159_2_n_34
    & sub_1159_2_n_17)));
 assign sub_1159_2_n_95 = ~(sub_1159_2_n_45 & (sub_1159_2_n_93 & (sub_1159_2_n_42 | sub_1159_2_n_5)));
 assign sub_1159_2_n_94 = ~(sub_1159_2_n_23 & (sub_1159_2_n_91 & (sub_1159_2_n_8 | sub_1159_2_n_13)));
 assign sub_1159_2_n_93 = ~(sub_1159_2_n_84 & sub_1159_2_n_64);
 assign sub_1159_2_n_92 = (sub_1159_2_n_88 | sub_1159_2_n_89);
 assign sub_1159_2_n_91 = ~(sub_1159_2_n_81 & sub_1159_2_n_77);
 assign sub_1159_2_n_87 = ~(sub_1159_2_n_43 | ~(sub_1159_2_n_31 | sub_1159_2_n_25));
 assign sub_1159_2_n_86 = ~(sub_1159_2_n_21 & (sub_1159_2_n_38 | sub_1159_2_n_28));
 assign sub_1159_2_n_90 = (sub_1159_2_n_76 & sub_1159_2_n_79);
 assign sub_1159_2_n_89 = ~(sub_1159_2_n_63 & sub_1159_2_n_77);
 assign sub_1159_2_n_88 = ~(sub_1159_2_n_75 & ~sub_1159_2_n_80);
 assign sub_1159_2_n_85 = ~(sub_1159_2_n_47 | ~(sub_1159_2_n_39 | sub_1159_2_n_9));
 assign sub_1159_2_n_84 = ~(sub_1159_2_n_24 & (sub_1159_2_n_27 | sub_1159_2_n_26));
 assign sub_1159_2_n_83 = ~(sub_1159_2_n_46 & (sub_1159_2_n_32 | sub_1159_2_n_40));
 assign sub_1159_2_n_82 = ~(sub_1159_2_n_20 & (sub_1159_2_n_6 | sub_1159_2_n_15));
 assign sub_1159_2_n_81 = ~(sub_1159_2_n_19 & (sub_1159_2_n_3 | sub_1159_2_n_14));
 assign sub_1159_2_n_74 = ~(sub_1159_2_n_17 & ~sub_1159_2_n_22);
 assign sub_1159_2_n_80 = (sub_1159_2_n_37 | sub_1159_2_n_15);
 assign sub_1159_2_n_73 = ~(sub_1159_2_n_7 & ~sub_1159_2_n_30);
 assign sub_1159_2_n_79 = ~(sub_1159_2_n_16 | sub_1159_2_n_28);
 assign sub_1159_2_n_78 = (sub_1159_2_n_36 | sub_1159_2_n_25);
 assign sub_1159_2_n_72 = ~(sub_1159_2_n_23 & ~sub_1159_2_n_13);
 assign sub_1159_2_n_71 = ~(sub_1159_2_n_24 & ~sub_1159_2_n_26);
 assign sub_1159_2_n_70 = ~(sub_1159_2_n_4 | ~sub_1159_2_n_39);
 assign sub_1159_2_n_77 = ~(sub_1159_2_n_29 | sub_1159_2_n_13);
 assign sub_1159_2_n_69 = (sub_1159_2_n_47 | sub_1159_2_n_9);
 assign sub_1159_2_n_68 = ~(sub_1159_2_n_29 | ~sub_1159_2_n_8);
 assign sub_1159_2_n_67 = ~(sub_1159_2_n_19 & ~sub_1159_2_n_14);
 assign sub_1159_2_n_76 = ~(sub_1159_2_n_40 | ~sub_1159_2_n_12);
 assign sub_1159_2_n_75 = ~(sub_1159_2_n_41 | ~sub_1159_2_n_17);
 assign sub_1159_2_n_66 = ~(sub_1159_2_n_3 & sub_1159_2_n_33);
 assign sub_1159_2_n_65 = ~(sub_1159_2_n_18 | ~sub_1159_2_n_42);
 assign sub_1159_2_n_61 = (sub_1159_2_n_7 & sub_1159_2_n_11);
 assign in1_139_0_ = ~(sub_1159_2_n_2 & ~(sub_1159_2_n_0 & n_1471));
 assign sub_1159_2_n_59 = ~(sub_1159_2_n_36 | ~sub_1159_2_n_31);
 assign sub_1159_2_n_58 = ~(sub_1159_2_n_37 | ~sub_1159_2_n_6);
 assign sub_1159_2_n_57 = (sub_1159_2_n_43 | sub_1159_2_n_25);
 assign sub_1159_2_n_56 = ~(sub_1159_2_n_34 | sub_1159_2_n_41);
 assign sub_1159_2_n_55 = ~(sub_1159_2_n_44 | ~sub_1159_2_n_11);
 assign sub_1159_2_n_64 = ~(sub_1159_2_n_18 | sub_1159_2_n_5);
 assign sub_1159_2_n_63 = ~(sub_1159_2_n_14 | ~sub_1159_2_n_33);
 assign sub_1159_2_n_54 = ~(sub_1159_2_n_16 | ~sub_1159_2_n_38);
 assign sub_1159_2_n_53 = ~(sub_1159_2_n_46 & ~sub_1159_2_n_40);
 assign sub_1159_2_n_52 = ~(sub_1159_2_n_32 & sub_1159_2_n_12);
 assign sub_1159_2_n_51 = ~(sub_1159_2_n_27 & sub_1159_2_n_10);
 assign sub_1159_2_n_50 = ~(sub_1159_2_n_45 & ~sub_1159_2_n_5);
 assign sub_1159_2_n_49 = ~(sub_1159_2_n_21 & ~sub_1159_2_n_28);
 assign sub_1159_2_n_62 = ~(sub_1159_2_n_26 | ~sub_1159_2_n_10);
 assign sub_1159_2_n_48 = ~(sub_1159_2_n_20 & ~sub_1159_2_n_15);
 assign sub_1159_2_n_35 = ~sub_1159_2_n_34;
 assign sub_1159_2_n_47 = ~(n_1570 | ~in1_137_4_);
 assign sub_1159_2_n_46 = ~(in1_137_12_ & ~n_1582);
 assign sub_1159_2_n_45 = ~(in1_137_10_ & ~n_1556);
 assign sub_1159_2_n_44 = ~(n_1580 | ~in1_137_2_);
 assign sub_1159_2_n_43 = ~(n_1528 | ~in1_137_6_);
 assign sub_1159_2_n_42 = ~(in1_137_9_ & ~n_1552);
 assign sub_1159_2_n_41 = ~(in1_137_17_ | ~n_1473);
 assign sub_1159_2_n_40 = ~(in1_137_12_ | ~n_1582);
 assign sub_1159_2_n_39 = ~(in1_137_3_ & ~n_1536);
 assign sub_1159_2_n_38 = ~(in1_137_13_ & ~n_1578);
 assign sub_1159_2_n_37 = ~(in1_137_15_ | ~n_1550);
 assign sub_1159_2_n_36 = ~(in1_137_5_ | ~n_1568);
 assign sub_1159_2_n_34 = ~(n_1473 | ~in1_137_17_);
 assign sub_1159_2_n_33 = ~(n_1566 & ~in1_137_19_);
 assign sub_1159_2_n_32 = ~(in1_137_11_ & ~n_1596);
 assign sub_1159_2_n_31 = ~(in1_137_5_ & ~n_1568);
 assign sub_1159_2_n_30 = ~(n_1478 | ~in1_137_1_);
 assign sub_1159_2_n_29 = ~(in1_137_21_ | ~n_1592);
 assign sub_1159_2_n_28 = ~(in1_137_14_ | ~n_1496);
 assign sub_1159_2_n_27 = ~(in1_137_7_ & ~n_1480);
 assign sub_1159_2_n_26 = ~(in1_137_8_ | ~n_1590);
 assign sub_1159_2_n_25 = ~(in1_137_6_ | ~n_1528);
 assign sub_1159_2_n_24 = ~(in1_137_8_ & ~n_1590);
 assign sub_1159_2_n_23 = ~(in1_137_22_ & ~n_1404);
 assign sub_1159_2_n_22 = ~(n_1559 | ~in1_137_18_);
 assign sub_1159_2_n_21 = ~(in1_137_14_ & ~n_1496);
 assign sub_1159_2_n_20 = ~(in1_137_16_ & ~n_1563);
 assign sub_1159_2_n_19 = ~(in1_137_20_ & ~n_1594);
 assign sub_1159_2_n_18 = ~(in1_137_9_ | ~n_1552);
 assign sub_1159_2_n_17 = ~(n_1559 & ~in1_137_18_);
 assign sub_1159_2_n_16 = ~(in1_137_13_ | ~n_1578);
 assign sub_1159_2_n_15 = ~(in1_137_16_ | ~n_1563);
 assign sub_1159_2_n_14 = ~(in1_137_20_ | ~n_1594);
 assign sub_1159_2_n_13 = ~(in1_137_22_ | ~n_1404);
 assign sub_1159_2_n_12 = ~(n_1596 & ~in1_137_11_);
 assign sub_1159_2_n_11 = ~(n_1580 & ~in1_137_2_);
 assign sub_1159_2_n_10 = ~(n_1480 & ~in1_137_7_);
 assign sub_1159_2_n_9 = ~(in1_137_4_ | ~n_1570);
 assign sub_1159_2_n_8 = ~(in1_137_21_ & ~n_1592);
 assign sub_1159_2_n_7 = ~(n_1478 & ~in1_137_1_);
 assign sub_1159_2_n_6 = ~(in1_137_15_ & ~n_1550);
 assign sub_1159_2_n_5 = ~(in1_137_10_ | ~n_1556);
 assign sub_1159_2_n_4 = ~(in1_137_3_ | ~n_1536);
 assign sub_1159_2_n_3 = ~(in1_137_19_ & ~n_1566);
 assign sub_1159_2_n_2 = ~(n_1544 & ~n_1471);
 assign sub_1159_2_n_1 = ~n_1587;
 assign sub_1159_2_n_0 = ~n_1544;
 assign in1_142_23_ = ~(sub_1180_2_n_148 ^ sub_1180_2_n_72);
 assign sub_1180_2_n_148 = ~(sub_1180_2_n_8 & (sub_1180_2_n_143 | sub_1180_2_n_29));
 assign in1_142_22_ = ~(sub_1180_2_n_143 ^ sub_1180_2_n_68);
 assign in1_142_21_ = ~(sub_1180_2_n_142 ^ sub_1180_2_n_67);
 assign in1_142_19_ = ~(sub_1180_2_n_141 ^ sub_1180_2_n_74);
 assign in1_142_15_ = ~(sub_1180_2_n_137 ^ sub_1180_2_n_49);
 assign sub_1180_2_n_143 = ~(sub_1180_2_n_82 | (sub_1180_2_n_132 & sub_1180_2_n_63));
 assign sub_1180_2_n_142 = ~(sub_1180_2_n_3 & ~(sub_1180_2_n_132 & sub_1180_2_n_33));
 assign sub_1180_2_n_141 = ~(sub_1180_2_n_35 & (sub_1180_2_n_131 | sub_1180_2_n_41));
 assign in1_142_20_ = ~(sub_1180_2_n_132 ^ sub_1180_2_n_66);
 assign in1_142_18_ = ~(sub_1180_2_n_131 ^ sub_1180_2_n_48);
 assign in1_142_17_ = ~(sub_1180_2_n_130 ^ sub_1180_2_n_59);
 assign sub_1180_2_n_137 = ~(sub_1180_2_n_38 & (sub_1180_2_n_127 | sub_1180_2_n_16));
 assign in1_142_24_ = ~(sub_1180_2_n_128 ^ in1_140_23_);
 assign in1_142_14_ = ~(sub_1180_2_n_127 ^ sub_1180_2_n_54);
 assign in1_142_13_ = ~(sub_1180_2_n_126 ^ sub_1180_2_n_53);
 assign in1_142_11_ = ~(sub_1180_2_n_125 ^ sub_1180_2_n_50);
 assign sub_1180_2_n_132 = ~(sub_1180_2_n_97 & (sub_1180_2_n_121 | sub_1180_2_n_89));
 assign sub_1180_2_n_131 = ~(sub_1180_2_n_83 | ~(sub_1180_2_n_121 | sub_1180_2_n_80));
 assign sub_1180_2_n_130 = ~(sub_1180_2_n_6 & (sub_1180_2_n_121 | sub_1180_2_n_37));
 assign in1_142_16_ = ~(sub_1180_2_n_121 ^ sub_1180_2_n_57);
 assign sub_1180_2_n_128 = ~(sub_1180_2_n_100 & ((sub_1180_2_n_101 | sub_1180_2_n_93) & (sub_1180_2_n_119
    | sub_1180_2_n_93)));
 assign sub_1180_2_n_127 = ~(sub_1180_2_n_84 | (sub_1180_2_n_118 & sub_1180_2_n_76));
 assign sub_1180_2_n_126 = ~(sub_1180_2_n_32 & ~(sub_1180_2_n_118 & sub_1180_2_n_12));
 assign sub_1180_2_n_125 = ~(sub_1180_2_n_42 & (sub_1180_2_n_117 | sub_1180_2_n_18));
 assign in1_142_12_ = ~(sub_1180_2_n_118 ^ sub_1180_2_n_52);
 assign in1_142_10_ = ~(sub_1180_2_n_117 ^ sub_1180_2_n_65);
 assign in1_142_9_ = ~(sub_1180_2_n_116 ^ sub_1180_2_n_71);
 assign sub_1180_2_n_121 = (sub_1180_2_n_119 & sub_1180_2_n_101);
 assign in1_142_7_ = ~(sub_1180_2_n_114 ^ sub_1180_2_n_56);
 assign sub_1180_2_n_119 = ~(sub_1180_2_n_113 & sub_1180_2_n_91);
 assign sub_1180_2_n_118 = (sub_1180_2_n_113 | sub_1180_2_n_96);
 assign sub_1180_2_n_117 = ~(sub_1180_2_n_86 | (sub_1180_2_n_110 & sub_1180_2_n_62));
 assign sub_1180_2_n_116 = ~(sub_1180_2_n_27 & ~(sub_1180_2_n_110 & sub_1180_2_n_10));
 assign in1_142_8_ = ~(sub_1180_2_n_110 ^ sub_1180_2_n_51);
 assign sub_1180_2_n_114 = ~(sub_1180_2_n_31 | (sub_1180_2_n_109 & sub_1180_2_n_36));
 assign sub_1180_2_n_113 = (sub_1180_2_n_62 & (sub_1180_2_n_64 & sub_1180_2_n_110));
 assign in1_142_6_ = ~(sub_1180_2_n_109 ^ sub_1180_2_n_58);
 assign in1_142_5_ = ~(sub_1180_2_n_108 ^ sub_1180_2_n_69);
 assign sub_1180_2_n_110 = ~(sub_1180_2_n_88 & ((sub_1180_2_n_85 | sub_1180_2_n_78) & (sub_1180_2_n_105
    | sub_1180_2_n_78)));
 assign sub_1180_2_n_109 = ~(sub_1180_2_n_105 & sub_1180_2_n_85);
 assign sub_1180_2_n_108 = ~(sub_1180_2_n_39 & (sub_1180_2_n_102 | sub_1180_2_n_4));
 assign in1_142_4_ = ~(sub_1180_2_n_102 ^ sub_1180_2_n_70);
 assign in1_142_3_ = ~(sub_1180_2_n_104 ^ sub_1180_2_n_55);
 assign sub_1180_2_n_105 = (sub_1180_2_n_4 | (sub_1180_2_n_9 | sub_1180_2_n_102));
 assign sub_1180_2_n_104 = ~(sub_1180_2_n_30 & ~(sub_1180_2_n_99 & sub_1180_2_n_7));
 assign in1_142_2_ = ~(sub_1180_2_n_99 ^ sub_1180_2_n_73);
 assign sub_1180_2_n_102 = ~(sub_1180_2_n_81 | (sub_1180_2_n_7 & (sub_1180_2_n_11 & sub_1180_2_n_99)));
 assign sub_1180_2_n_101 = ~(sub_1180_2_n_87 | ((sub_1180_2_n_96 & sub_1180_2_n_91) | (sub_1180_2_n_84
    & sub_1180_2_n_79)));
 assign sub_1180_2_n_100 = ~(sub_1180_2_n_95 | ~(sub_1180_2_n_97 | sub_1180_2_n_90));
 assign sub_1180_2_n_99 = ((sub_1180_2_n_2 & in1_140_0_) | ((in1_140_0_ & sub_1180_2_n_1) | (sub_1180_2_n_1
    & sub_1180_2_n_2)));
 assign in1_142_1_ = (in1_140_0_ ^ (sub_1180_2_n_1 ^ sub_1180_2_n_2));
 assign sub_1180_2_n_97 = ~(sub_1180_2_n_22 | ((sub_1180_2_n_83 & sub_1180_2_n_75) | (sub_1180_2_n_34
    & sub_1180_2_n_17)));
 assign sub_1180_2_n_96 = ~(sub_1180_2_n_45 & (sub_1180_2_n_94 & (sub_1180_2_n_42 | sub_1180_2_n_5)));
 assign sub_1180_2_n_95 = ~(sub_1180_2_n_23 & (sub_1180_2_n_92 & (sub_1180_2_n_8 | sub_1180_2_n_13)));
 assign sub_1180_2_n_94 = ~(sub_1180_2_n_86 & sub_1180_2_n_64);
 assign sub_1180_2_n_93 = (sub_1180_2_n_89 | sub_1180_2_n_90);
 assign sub_1180_2_n_92 = ~(sub_1180_2_n_82 & sub_1180_2_n_77);
 assign sub_1180_2_n_88 = ~(sub_1180_2_n_43 | (sub_1180_2_n_31 & sub_1180_2_n_25));
 assign sub_1180_2_n_87 = ~(sub_1180_2_n_21 & (sub_1180_2_n_38 | sub_1180_2_n_28));
 assign sub_1180_2_n_91 = (sub_1180_2_n_76 & sub_1180_2_n_79);
 assign sub_1180_2_n_90 = ~(sub_1180_2_n_63 & sub_1180_2_n_77);
 assign sub_1180_2_n_89 = ~(sub_1180_2_n_75 & ~sub_1180_2_n_80);
 assign sub_1180_2_n_81 = ~(sub_1180_2_n_61 & sub_1180_2_n_44);
 assign sub_1180_2_n_86 = ~(sub_1180_2_n_24 & (sub_1180_2_n_27 | sub_1180_2_n_26));
 assign sub_1180_2_n_85 = ~(sub_1180_2_n_47 | ~(sub_1180_2_n_39 | sub_1180_2_n_9));
 assign sub_1180_2_n_84 = ~(sub_1180_2_n_46 & (sub_1180_2_n_32 | sub_1180_2_n_40));
 assign sub_1180_2_n_83 = ~(sub_1180_2_n_20 & (sub_1180_2_n_6 | sub_1180_2_n_15));
 assign sub_1180_2_n_82 = ~(sub_1180_2_n_19 & (sub_1180_2_n_3 | sub_1180_2_n_14));
 assign sub_1180_2_n_74 = ~(sub_1180_2_n_17 & ~sub_1180_2_n_22);
 assign sub_1180_2_n_80 = (sub_1180_2_n_37 | sub_1180_2_n_15);
 assign sub_1180_2_n_73 = ~(sub_1180_2_n_30 & sub_1180_2_n_7);
 assign sub_1180_2_n_79 = ~(sub_1180_2_n_16 | sub_1180_2_n_28);
 assign sub_1180_2_n_78 = ~(sub_1180_2_n_36 & sub_1180_2_n_25);
 assign sub_1180_2_n_72 = ~(sub_1180_2_n_23 & ~sub_1180_2_n_13);
 assign sub_1180_2_n_71 = ~(sub_1180_2_n_24 & ~sub_1180_2_n_26);
 assign sub_1180_2_n_70 = ~(sub_1180_2_n_4 | ~sub_1180_2_n_39);
 assign sub_1180_2_n_77 = ~(sub_1180_2_n_29 | sub_1180_2_n_13);
 assign sub_1180_2_n_69 = (sub_1180_2_n_47 | sub_1180_2_n_9);
 assign sub_1180_2_n_68 = ~(sub_1180_2_n_29 | ~sub_1180_2_n_8);
 assign sub_1180_2_n_67 = ~(sub_1180_2_n_19 & ~sub_1180_2_n_14);
 assign sub_1180_2_n_76 = ~(sub_1180_2_n_40 | ~sub_1180_2_n_12);
 assign sub_1180_2_n_75 = ~(sub_1180_2_n_41 | ~sub_1180_2_n_17);
 assign sub_1180_2_n_66 = ~(sub_1180_2_n_3 & sub_1180_2_n_33);
 assign sub_1180_2_n_65 = ~(sub_1180_2_n_18 | ~sub_1180_2_n_42);
 assign sub_1180_2_n_61 = ~(sub_1180_2_n_11 & ~sub_1180_2_n_30);
 assign in1_142_0_ = ~(sub_1180_2_n_2 & ~(sub_1180_2_n_0 & n_1400));
 assign sub_1180_2_n_59 = ~(sub_1180_2_n_20 & ~sub_1180_2_n_15);
 assign sub_1180_2_n_58 = ~(sub_1180_2_n_36 & ~sub_1180_2_n_31);
 assign sub_1180_2_n_57 = ~(sub_1180_2_n_37 | ~sub_1180_2_n_6);
 assign sub_1180_2_n_56 = ~(sub_1180_2_n_43 | ~sub_1180_2_n_25);
 assign sub_1180_2_n_55 = ~(sub_1180_2_n_44 & sub_1180_2_n_11);
 assign sub_1180_2_n_64 = ~(sub_1180_2_n_18 | sub_1180_2_n_5);
 assign sub_1180_2_n_63 = ~(sub_1180_2_n_14 | ~sub_1180_2_n_33);
 assign sub_1180_2_n_54 = ~(sub_1180_2_n_16 | ~sub_1180_2_n_38);
 assign sub_1180_2_n_53 = ~(sub_1180_2_n_46 & ~sub_1180_2_n_40);
 assign sub_1180_2_n_52 = ~(sub_1180_2_n_32 & sub_1180_2_n_12);
 assign sub_1180_2_n_51 = ~(sub_1180_2_n_27 & sub_1180_2_n_10);
 assign sub_1180_2_n_50 = ~(sub_1180_2_n_45 & ~sub_1180_2_n_5);
 assign sub_1180_2_n_49 = ~(sub_1180_2_n_21 & ~sub_1180_2_n_28);
 assign sub_1180_2_n_62 = ~(sub_1180_2_n_26 | ~sub_1180_2_n_10);
 assign sub_1180_2_n_48 = ~(sub_1180_2_n_34 | sub_1180_2_n_41);
 assign sub_1180_2_n_35 = ~sub_1180_2_n_34;
 assign sub_1180_2_n_47 = ~(n_1570 | ~in1_140_4_);
 assign sub_1180_2_n_46 = ~(in1_140_12_ & ~n_1582);
 assign sub_1180_2_n_45 = ~(in1_140_10_ & ~n_1556);
 assign sub_1180_2_n_44 = ~(in1_140_2_ & ~n_1580);
 assign sub_1180_2_n_43 = ~(n_1528 | ~in1_140_6_);
 assign sub_1180_2_n_42 = ~(in1_140_9_ & ~n_1552);
 assign sub_1180_2_n_41 = ~(in1_140_17_ | ~n_1473);
 assign sub_1180_2_n_40 = ~(in1_140_12_ | ~n_1582);
 assign sub_1180_2_n_39 = ~(in1_140_3_ & ~n_1536);
 assign sub_1180_2_n_38 = ~(in1_140_13_ & ~n_1578);
 assign sub_1180_2_n_37 = ~(in1_140_15_ | ~n_1550);
 assign sub_1180_2_n_36 = ~(n_1568 & ~in1_140_5_);
 assign sub_1180_2_n_34 = ~(n_1473 | ~in1_140_17_);
 assign sub_1180_2_n_33 = ~(n_1566 & ~in1_140_19_);
 assign sub_1180_2_n_32 = ~(in1_140_11_ & ~n_1596);
 assign sub_1180_2_n_31 = ~(n_1568 | ~in1_140_5_);
 assign sub_1180_2_n_30 = ~(in1_140_1_ & ~n_1478);
 assign sub_1180_2_n_29 = ~(in1_140_21_ | ~n_1592);
 assign sub_1180_2_n_28 = ~(in1_140_14_ | ~n_1496);
 assign sub_1180_2_n_27 = ~(in1_140_7_ & ~n_1480);
 assign sub_1180_2_n_26 = ~(in1_140_8_ | ~n_1590);
 assign sub_1180_2_n_25 = ~(n_1528 & ~in1_140_6_);
 assign sub_1180_2_n_24 = ~(in1_140_8_ & ~n_1590);
 assign sub_1180_2_n_23 = ~(in1_140_22_ & ~n_1404);
 assign sub_1180_2_n_22 = ~(n_1559 | ~in1_140_18_);
 assign sub_1180_2_n_21 = ~(in1_140_14_ & ~n_1496);
 assign sub_1180_2_n_20 = ~(in1_140_16_ & ~n_1563);
 assign sub_1180_2_n_19 = ~(in1_140_20_ & ~n_1594);
 assign sub_1180_2_n_18 = ~(in1_140_9_ | ~n_1552);
 assign sub_1180_2_n_17 = ~(n_1559 & ~in1_140_18_);
 assign sub_1180_2_n_16 = ~(in1_140_13_ | ~n_1578);
 assign sub_1180_2_n_15 = ~(in1_140_16_ | ~n_1563);
 assign sub_1180_2_n_14 = ~(in1_140_20_ | ~n_1594);
 assign sub_1180_2_n_13 = ~(in1_140_22_ | ~n_1404);
 assign sub_1180_2_n_12 = ~(n_1596 & ~in1_140_11_);
 assign sub_1180_2_n_11 = ~(n_1580 & ~in1_140_2_);
 assign sub_1180_2_n_10 = ~(n_1480 & ~in1_140_7_);
 assign sub_1180_2_n_9 = ~(in1_140_4_ | ~n_1570);
 assign sub_1180_2_n_8 = ~(in1_140_21_ & ~n_1592);
 assign sub_1180_2_n_7 = ~(n_1478 & ~in1_140_1_);
 assign sub_1180_2_n_6 = ~(in1_140_15_ & ~n_1550);
 assign sub_1180_2_n_5 = ~(in1_140_10_ | ~n_1556);
 assign sub_1180_2_n_4 = ~(in1_140_3_ | ~n_1536);
 assign sub_1180_2_n_3 = ~(in1_140_19_ & ~n_1566);
 assign sub_1180_2_n_2 = ~(n_1544 & ~n_1400);
 assign sub_1180_2_n_1 = ~n_1587;
 assign sub_1180_2_n_0 = ~n_1544;
 assign in1_145_24_ = ~(sub_1199_2_n_78 ^ in1_143_23_);
 assign sub_1199_2_n_78 = ~(sub_1199_2_n_77 & (sub_1199_2_n_76 & (sub_1199_2_n_74 | sub_1199_2_n_62)));
 assign sub_1199_2_n_77 = ~(sub_1199_2_n_73 & (sub_1199_2_n_55 & (sub_1199_2_n_75 | sub_1199_2_n_70)));
 assign sub_1199_2_n_76 = ~(sub_1199_2_n_60 | (sub_1199_2_n_71 | (sub_1199_2_n_59 & sub_1199_2_n_52)));
 assign sub_1199_2_n_75 = ~(sub_1199_2_n_33 | (sub_1199_2_n_43 | (sub_1199_2_n_53 | sub_1199_2_n_72)));
 assign sub_1199_2_n_74 = ~((sub_1199_2_n_1 & sub_1199_2_n_69) | (sub_1199_2_n_68 & sub_1199_2_n_0));
 assign sub_1199_2_n_73 = (sub_1199_2_n_67 & (sub_1199_2_n_52 & (sub_1199_2_n_39 & sub_1199_2_n_23)));
 assign sub_1199_2_n_72 = ~((sub_1199_2_n_22 & (sub_1199_2_n_29 & sub_1199_2_n_66)) | (sub_1199_2_n_45
    & sub_1199_2_n_29));
 assign sub_1199_2_n_71 = ~(sub_1199_2_n_62 | ((sub_1199_2_n_61 & sub_1199_2_n_32) | (sub_1199_2_n_57
    & sub_1199_2_n_48)));
 assign sub_1199_2_n_70 = ~(sub_1199_2_n_47 & (sub_1199_2_n_65 & (n_1528 | sub_1199_2_n_5)));
 assign sub_1199_2_n_69 = ~(sub_1199_2_n_51 & (sub_1199_2_n_64 & (n_1556 | sub_1199_2_n_6)));
 assign sub_1199_2_n_68 = ~(sub_1199_2_n_50 & ((n_1496 | sub_1199_2_n_13) & (sub_1199_2_n_58 | sub_1199_2_n_54)));
 assign sub_1199_2_n_67 = ~(sub_1199_2_n_26 | (sub_1199_2_n_54 | (sub_1199_2_n_21 | ~sub_1199_2_n_56)));
 assign sub_1199_2_n_66 = ~(sub_1199_2_n_63 & (sub_1199_2_n_36 | n_1587));
 assign sub_1199_2_n_65 = (sub_1199_2_n_46 | (sub_1199_2_n_43 | sub_1199_2_n_53));
 assign sub_1199_2_n_64 = ~(sub_1199_2_n_44 & (sub_1199_2_n_39 & (sub_1199_2_n_40 & sub_1199_2_n_35)));
 assign sub_1199_2_n_63 = ~(in1_143_0_ & ~(sub_1199_2_n_36 & n_1587));
 assign sub_1199_2_n_62 = ~(sub_1199_2_n_38 & (sub_1199_2_n_23 & sub_1199_2_n_52));
 assign sub_1199_2_n_61 = ~(sub_1199_2_n_30 & (sub_1199_2_n_25 | sub_1199_2_n_28));
 assign sub_1199_2_n_60 = ~((n_1592 | (sub_1199_2_n_11 | sub_1199_2_n_42)) & (n_1404 | sub_1199_2_n_10));
 assign sub_1199_2_n_59 = ~(sub_1199_2_n_49 & ~(sub_1199_2_n_17 & in1_143_20_));
 assign sub_1199_2_n_58 = ~((sub_1199_2_n_4 & (in1_143_11_ & sub_1199_2_n_27)) | (sub_1199_2_n_12 & in1_143_12_));
 assign sub_1199_2_n_57 = ~(sub_1199_2_n_31 | (sub_1199_2_n_28 | (sub_1199_2_n_14 & in1_143_16_)));
 assign sub_1199_2_n_56 = (sub_1199_2_n_30 & (sub_1199_2_n_37 & (sub_1199_2_n_25 & sub_1199_2_n_34)));
 assign sub_1199_2_n_55 = (sub_1199_2_n_20 & (sub_1199_2_n_40 & (sub_1199_2_n_35 & sub_1199_2_n_38)));
 assign sub_1199_2_n_51 = ~(in1_143_9_ & (sub_1199_2_n_35 & ~n_1552));
 assign sub_1199_2_n_50 = ~(in1_143_13_ & (sub_1199_2_n_24 & ~n_1578));
 assign sub_1199_2_n_54 = ~(sub_1199_2_n_24 & ~(sub_1199_2_n_8 & n_1578));
 assign sub_1199_2_n_53 = ~(sub_1199_2_n_41 & ~(sub_1199_2_n_19 & n_1568));
 assign sub_1199_2_n_52 = ~(sub_1199_2_n_42 | (sub_1199_2_n_11 & n_1592));
 assign sub_1199_2_n_49 = ~(in1_143_19_ & (sub_1199_2_n_23 & ~n_1566));
 assign sub_1199_2_n_48 = ~(in1_143_15_ & (sub_1199_2_n_37 & ~n_1550));
 assign sub_1199_2_n_47 = ~(in1_143_5_ & (sub_1199_2_n_41 & ~n_1568));
 assign sub_1199_2_n_46 = ~((sub_1199_2_n_3 & in1_143_3_) | (sub_1199_2_n_7 & in1_143_4_));
 assign sub_1199_2_n_45 = ~((n_1478 | sub_1199_2_n_18) & (n_1580 | sub_1199_2_n_16));
 assign sub_1199_2_n_44 = ~((n_1480 | sub_1199_2_n_15) & (n_1590 | sub_1199_2_n_9));
 assign sub_1199_2_n_34 = ~(n_1550 & ~in1_143_15_);
 assign sub_1199_2_n_33 = ~(in1_143_3_ | sub_1199_2_n_3);
 assign sub_1199_2_n_43 = ~(in1_143_4_ | sub_1199_2_n_7);
 assign sub_1199_2_n_42 = ~(in1_143_22_ | ~n_1404);
 assign sub_1199_2_n_41 = ~(sub_1199_2_n_5 & n_1528);
 assign sub_1199_2_n_40 = ~(n_1552 & ~in1_143_9_);
 assign sub_1199_2_n_39 = ~(sub_1199_2_n_9 & n_1590);
 assign sub_1199_2_n_38 = ~(n_1566 & ~in1_143_19_);
 assign sub_1199_2_n_37 = (in1_143_16_ | sub_1199_2_n_14);
 assign sub_1199_2_n_36 = ~(n_1398 | ~n_1544);
 assign sub_1199_2_n_35 = ~(sub_1199_2_n_6 & n_1556);
 assign sub_1199_2_n_32 = ~sub_1199_2_n_31;
 assign sub_1199_2_n_27 = ~sub_1199_2_n_26;
 assign sub_1199_2_n_22 = ~(sub_1199_2_n_18 & n_1478);
 assign sub_1199_2_n_21 = ~(in1_143_11_ | sub_1199_2_n_4);
 assign sub_1199_2_n_20 = ~(sub_1199_2_n_15 & n_1480);
 assign sub_1199_2_n_31 = ~(n_1559 | ~in1_143_18_);
 assign sub_1199_2_n_30 = ~(n_1559 & ~in1_143_18_);
 assign sub_1199_2_n_29 = ~(sub_1199_2_n_16 & n_1580);
 assign sub_1199_2_n_28 = ~(n_1473 | ~in1_143_17_);
 assign sub_1199_2_n_26 = ~(in1_143_12_ | sub_1199_2_n_12);
 assign sub_1199_2_n_25 = ~(n_1473 & ~in1_143_17_);
 assign sub_1199_2_n_24 = ~(sub_1199_2_n_13 & n_1496);
 assign sub_1199_2_n_23 = (in1_143_20_ | sub_1199_2_n_17);
 assign sub_1199_2_n_19 = ~in1_143_5_;
 assign sub_1199_2_n_18 = ~in1_143_1_;
 assign sub_1199_2_n_17 = ~n_1594;
 assign sub_1199_2_n_16 = ~in1_143_2_;
 assign sub_1199_2_n_15 = ~in1_143_7_;
 assign sub_1199_2_n_14 = ~n_1563;
 assign sub_1199_2_n_13 = ~in1_143_14_;
 assign sub_1199_2_n_12 = ~n_1582;
 assign sub_1199_2_n_11 = ~in1_143_21_;
 assign sub_1199_2_n_10 = ~in1_143_22_;
 assign sub_1199_2_n_9 = ~in1_143_8_;
 assign sub_1199_2_n_8 = ~in1_143_13_;
 assign sub_1199_2_n_7 = ~n_1570;
 assign sub_1199_2_n_6 = ~in1_143_10_;
 assign sub_1199_2_n_5 = ~in1_143_6_;
 assign sub_1199_2_n_4 = ~n_1596;
 assign sub_1199_2_n_3 = ~n_1536;
 assign sub_1199_2_n_1 = sub_1199_2_n_67;
 assign sub_1199_2_n_0 = sub_1199_2_n_56;
endmodule

